//The Netlist from Uncle 
module ncl_up_counter ( t_out  ,  f_out  ,  t_enable  ,  f_enable  ,  t_clr  ,  f_clr  ,  reset  ,  ackout  ,  ackin );
  input ackin ;
  output ackout ;
  input reset ;
  input f_clr ;
  input t_clr ;
  input f_enable ;
  input t_enable ;
  output [7:0] f_out ;
  output [7:0] t_out ;

  wire [7:0] f_next_out ;
  wire [7:0] t_next_out ;
  wire [7:0] f_out_now ;
  wire [7:0] t_out_now ;
  wire n1_N_15 ;
  wire ki_N_0 ;
  wire ki_N ;
  wire acknet13 ;
  wire acknet12 ;
  wire acknet11 ;
  wire acknet10 ;
  wire acknet9 ;
  wire acknet8 ;
  wire acknet7 ;
  wire acknet6 ;
  wire acknet5 ;
  wire acknet4 ;
  wire acknet3 ;
  wire acknet2 ;
  wire s0_start ;
  wire s1_start ;
  wire s1_done ;
  wire f_n2 ;
  wire t_n2 ;
  wire f_n1 ;
  wire t_n1 ;
  wire f_n6 ;
  wire t_n6 ;
  wire f_n5 ;
  wire t_n5 ;
  wire f_n8 ;
  wire t_n8 ;
  wire f_n7 ;
  wire t_n7 ;
  wire f_n10 ;
  wire t_n10 ;
  wire f_n9 ;
  wire t_n9 ;
  wire f_n12 ;
  wire t_n12 ;
  wire f_n11 ;
  wire t_n11 ;
  wire f_n14 ;
  wire t_n14 ;
  wire f_n13 ;
  wire t_n13 ;
  wire f_n16 ;
  wire t_n16 ;
  wire f_n15 ;
  wire t_n15 ;
  wire f_n18 ;
  wire t_n18 ;
  wire f_n3 ;
  wire t_n3 ;
  wire f_n17 ;
  wire t_n17 ;
  wire f_n4 ;
  wire t_n4 ;
  wire f_n19 ;
  wire t_n19 ;
  wire f_n20 ;
  wire t_n20 ;
  wire \f_dout_master/genblk1[0].g0/n1 ;
  wire \t_dout_master/genblk1[0].g0/n1 ;
  wire \f_dout_slave/genblk1[7].g0/n1 ;
  wire \t_dout_slave/genblk1[7].g0/n1 ;
  wire \f_dout_slave/genblk1[6].g0/n1 ;
  wire \t_dout_slave/genblk1[6].g0/n1 ;
  wire \f_dout_slave/genblk1[5].g0/n1 ;
  wire \t_dout_slave/genblk1[5].g0/n1 ;
  wire \f_dout_slave/genblk1[4].g0/n1 ;
  wire \t_dout_slave/genblk1[4].g0/n1 ;
  wire \f_dout_slave/genblk1[3].g0/n1 ;
  wire \t_dout_slave/genblk1[3].g0/n1 ;
  wire \f_dout_slave/genblk1[2].g0/n1 ;
  wire \t_dout_slave/genblk1[2].g0/n1 ;
  wire \f_dout_slave/genblk1[1].g0/n1 ;
  wire \t_dout_slave/genblk1[1].g0/n1 ;
  wire \f_dout_slave/genblk1[0].g0/n1 ;
  wire \t_dout_slave/genblk1[0].g0/n1 ;
  wire \f_dout_master/genblk1[7].g0/n1 ;
  wire \t_dout_master/genblk1[7].g0/n1 ;
  wire \f_dout_master/genblk1[6].g0/n1 ;
  wire \t_dout_master/genblk1[6].g0/n1 ;
  wire \f_dout_master/genblk1[5].g0/n1 ;
  wire \t_dout_master/genblk1[5].g0/n1 ;
  wire \f_dout_master/genblk1[4].g0/n1 ;
  wire \t_dout_master/genblk1[4].g0/n1 ;
  wire \f_dout_master/genblk1[3].g0/n1 ;
  wire \t_dout_master/genblk1[3].g0/n1 ;
  wire \f_dout_master/genblk1[2].g0/n1 ;
  wire \t_dout_master/genblk1[2].g0/n1 ;
  wire s1 ;
  wire \f_dout_master/genblk1[1].g0/n1 ;
  wire \t_dout_master/genblk1[1].g0/n1 ;
  wire f_N5 ;
  wire t_N5 ;
  wire f_N6 ;
  wire t_N6 ;
  wire f_N7 ;
  wire t_N7 ;
  wire f_n21 ;
  wire t_n21 ;
  wire f_N8 ;
  wire t_N8 ;
  wire f_n22 ;
  wire t_n22 ;
  wire f_N9 ;
  wire t_N9 ;
  wire f_n23 ;
  wire t_n23 ;
  wire f_N10 ;
  wire t_N10 ;
  wire f_n24 ;
  wire t_n24 ;
  wire f_N11 ;
  wire t_N11 ;
  wire f_n25 ;
  wire t_n25 ;
  wire f_n26 ;
  wire t_n26 ;
  wire f_N12 ;
  wire t_N12 ;
  wire s0 ;
  wire n1_N ;
  wire n1_N_0 ;
  wire n1_N_1 ;
  wire n1_N_2 ;
  wire n1_N_3 ;
  wire n1_N_4 ;
  wire n1_N_5 ;
  wire n1_N_6 ;
  wire n1_N_7 ;
  wire n1_N_8 ;
  wire n1_N_9 ;
  wire n1_N_10 ;
  wire n1_N_11 ;
  wire n1_N_12 ;
  wire n1_N_13 ;
  wire n1_N_14 ;
  wire en_b_N ;
  wire t_enable ;
  wire f_enable ;
  wire t_clr ;
  wire f_clr ;
  wire reset ;
  wire ackout ;
  wire ackin ;
  assign s1_done = ki_N_0 ; 
  assign t_n20 = f_enable ; 
  assign ackout = acknet13 ; 
  assign t_n19 = f_clr ; 
  assign s1 = s1_start ; 
  assign f_N5 = t_out_now[0] ; 
  assign f_n20 = t_enable ; 
  assign f_n19 = t_clr ; 
  assign t_N5 = f_out_now[0] ; 
  and2x4  u1_U_U_1 (.a ( n1_N_15 ) , .b ( s0_start ) , .y ( s0 ));
  nor2  u1_U_U_0 (.a ( ki_N ) , .b ( n1_N_15 ) , .y ( s1_start ));
  nc2p  u1_U_U (.a ( s0_start ) , .b ( ki_N ) , .y ( n1_N_15 ));
  inv  u2_U_0 (.a ( acknet12 ) , .y ( ki_N_0 ));
  inv  u1_U_0 (.a ( acknet9 ) , .y ( ki_N ));
  th22  cgate11 (.a ( acknet6 ) , .b ( acknet6 ) , .y ( acknet13 ));
  th33  cgate10 (.a ( n1_N_6 ) , .b ( acknet11 ) , .c ( acknet10 ) , .y ( acknet12 ));
  th44  cgate9 (.a ( n1_N_7 ) , .b ( n1_N_9 ) , .c ( n1_N_11 ) , .d ( n1_N_13 ) , .y ( acknet11 ));
  th44  cgate8 (.a ( n1_N_8 ) , .b ( n1_N_10 ) , .c ( n1_N_12 ) , .d ( ackin ) , .y ( acknet10 ));
  th22  cgate7 (.a ( acknet8 ) , .b ( acknet7 ) , .y ( acknet9 ));
  th44  cgate6 (.a ( n1_N_5 ) , .b ( n1_N_0 ) , .c ( n1_N_2 ) , .d ( n1_N_4 ) , .y ( acknet8 ));
  th44  cgate5 (.a ( n1_N_14 ) , .b ( n1_N ) , .c ( n1_N_1 ) , .d ( n1_N_3 ) , .y ( acknet7 ));
  th44  cgate4 (.a ( acknet5 ) , .b ( acknet4 ) , .c ( acknet3 ) , .d ( acknet2 ) , .y ( acknet6 ));
  th33r  cgate3 (.a ( s0 ) , .b ( n1_N ) , .c ( n1_N_14 ) , .rsb ( reset ) , .y ( acknet5 ));
  th33r  cgate2 (.a ( s0 ) , .b ( n1_N_1 ) , .c ( n1_N_0 ) , .rsb ( reset ) , .y ( acknet4 ));
  th33r  cgate1 (.a ( s0 ) , .b ( n1_N_3 ) , .c ( n1_N_2 ) , .rsb ( reset ) , .y ( acknet3 ));
  th33r  cgate0 (.a ( s0 ) , .b ( n1_N_5 ) , .c ( n1_N_4 ) , .rsb ( reset ) , .y ( acknet2 ));
  th24comp  U45_U (.y ( t_N12 ) , .d ( f_out_now[7] ) , .c ( f_n26 ) , .b ( t_n26 ) , .a ( t_out_now[7] ));
  th24comp  U45_U_0 (.y ( f_N12 ) , .d ( f_out_now[7] ) , .c ( t_n26 ) , .b ( f_n26 ) , .a ( t_out_now[7] ));
  thand0  U44_U (.y ( f_n26 ) , .d ( t_n25 ) , .c ( t_out_now[6] ) , .b ( f_n25 ) , .a ( f_out_now[6] ));
  th22  U44_U_0 (.y ( t_n26 ) , .b ( t_n25 ) , .a ( t_out_now[6] ));
  th24comp  U43_U (.y ( t_N11 ) , .d ( f_out_now[6] ) , .c ( f_n25 ) , .b ( t_n25 ) , .a ( t_out_now[6] ));
  th24comp  U43_U_0 (.y ( f_N11 ) , .d ( f_out_now[6] ) , .c ( t_n25 ) , .b ( f_n25 ) , .a ( t_out_now[6] ));
  thand0  U42_U (.y ( f_n25 ) , .d ( t_out_now[5] ) , .c ( t_n24 ) , .b ( f_out_now[5] ) , .a ( f_n24 ));
  th22  U42_U_0 (.y ( t_n25 ) , .b ( t_out_now[5] ) , .a ( t_n24 ));
  th24comp  U41_U (.y ( t_N10 ) , .d ( f_out_now[5] ) , .c ( f_n24 ) , .b ( t_n24 ) , .a ( t_out_now[5] ));
  th24comp  U41_U_0 (.y ( f_N10 ) , .d ( f_out_now[5] ) , .c ( t_n24 ) , .b ( f_n24 ) , .a ( t_out_now[5] ));
  thand0  U40_U (.y ( f_n24 ) , .d ( t_n23 ) , .c ( t_out_now[4] ) , .b ( f_n23 ) , .a ( f_out_now[4] ));
  th22  U40_U_0 (.y ( t_n24 ) , .b ( t_n23 ) , .a ( t_out_now[4] ));
  th24comp  U39_U (.y ( t_N9 ) , .d ( f_out_now[4] ) , .c ( f_n23 ) , .b ( t_n23 ) , .a ( t_out_now[4] ));
  th24comp  U39_U_0 (.y ( f_N9 ) , .d ( f_out_now[4] ) , .c ( t_n23 ) , .b ( f_n23 ) , .a ( t_out_now[4] ));
  thand0  U38_U (.y ( f_n23 ) , .d ( t_n22 ) , .c ( t_out_now[3] ) , .b ( f_n22 ) , .a ( f_out_now[3] ));
  th22  U38_U_0 (.y ( t_n23 ) , .b ( t_n22 ) , .a ( t_out_now[3] ));
  th24comp  U37_U (.y ( t_N8 ) , .d ( f_out_now[3] ) , .c ( f_n22 ) , .b ( t_n22 ) , .a ( t_out_now[3] ));
  th24comp  U37_U_0 (.y ( f_N8 ) , .d ( f_out_now[3] ) , .c ( t_n22 ) , .b ( f_n22 ) , .a ( t_out_now[3] ));
  thand0  U36_U (.y ( f_n22 ) , .d ( t_n21 ) , .c ( t_out_now[2] ) , .b ( f_n21 ) , .a ( f_out_now[2] ));
  th22  U36_U_0 (.y ( t_n22 ) , .b ( t_n21 ) , .a ( t_out_now[2] ));
  th24comp  U35_U (.y ( t_N7 ) , .d ( f_out_now[2] ) , .c ( f_n21 ) , .b ( t_n21 ) , .a ( t_out_now[2] ));
  th24comp  U35_U_0 (.y ( f_N7 ) , .d ( f_out_now[2] ) , .c ( t_n21 ) , .b ( f_n21 ) , .a ( t_out_now[2] ));
  thand0  U34_U (.y ( f_n21 ) , .d ( t_out_now[0] ) , .c ( t_out_now[1] ) , .b ( f_out_now[0] ) , .a ( f_out_now[1] ));
  th22  U34_U_0 (.y ( t_n21 ) , .b ( t_out_now[0] ) , .a ( t_out_now[1] ));
  th24comp  U33_U (.y ( t_N6 ) , .d ( f_out_now[1] ) , .c ( f_out_now[0] ) , .b ( t_out_now[0] ) , .a ( t_out_now[1] ));
  th24comp  U33_U_0 (.y ( f_N6 ) , .d ( f_out_now[1] ) , .c ( t_out_now[0] ) , .b ( f_out_now[0] ) , .a ( t_out_now[1] ));
  srdreg  \dout_master/genblk1[1].g0/g0_U (.ackout ( n1_N ) , 
  
  .f_q ( \f_dout_master/genblk1[1].g0/n1 )
  
   , .t_q ( \t_dout_master/genblk1[1].g0/n1 ) , .f_d ( f_next_out[1] ) , .t_d ( t_next_out[1] ));
  and2  \dout_master/genblk1[1].g0/g1_U (.y ( t_out[1] ) , .b ( s1_start ) , .a ( \t_dout_master/genblk1[1].g0/n1 ));
  and2  \dout_master/genblk1_1_.g0/g1_U_0 (.y ( f_out[1] ) , .b ( s1_start ) , .a ( \f_dout_master/genblk1[1].g0/n1 ));
  srdreg  \dout_master/genblk1[2].g0/g0_U (.ackout ( n1_N_0 ) , .f_q ( \f_dout_master/genblk1[2].g0/n1 ) , .t_q ( \t_dout_master/genblk1[2].g0/n1 ) , .f_d ( f_next_out[2] ) , .t_d ( t_next_out[2] ));
  and2  \dout_master/genblk1[2].g0/g1_U (.y ( t_out[2] ) , .b ( s1_start ) , .a ( \t_dout_master/genblk1[2].g0/n1 ));
  and2  \dout_master/genblk1_2_.g0/g1_U_0 (.y ( f_out[2] ) , .b ( s1_start ) , .a ( \f_dout_master/genblk1[2].g0/n1 ));
  srdreg  \dout_master/genblk1[3].g0/g0_U (.ackout ( n1_N_1 ) , .f_q ( \f_dout_master/genblk1[3].g0/n1 ) , .t_q ( \t_dout_master/genblk1[3].g0/n1 ) , .f_d ( f_next_out[3] ) , .t_d ( t_next_out[3] ));
  and2  \dout_master/genblk1[3].g0/g1_U (.y ( t_out[3] ) , .b ( s1_start ) , .a ( \t_dout_master/genblk1[3].g0/n1 ));
  and2  \dout_master/genblk1_3_.g0/g1_U_0 (.y ( f_out[3] ) , .b ( s1_start ) , .a ( \f_dout_master/genblk1[3].g0/n1 ));
  srdreg  \dout_master/genblk1[4].g0/g0_U (.ackout ( n1_N_2 ) , .f_q ( \f_dout_master/genblk1[4].g0/n1 ) , .t_q ( \t_dout_master/genblk1[4].g0/n1 ) , .f_d ( f_next_out[4] ) , .t_d ( t_next_out[4] ));
  and2  \dout_master/genblk1[4].g0/g1_U (.y ( t_out[4] ) , .b ( s1_start ) , .a ( \t_dout_master/genblk1[4].g0/n1 ));
  and2  \dout_master/genblk1_4_.g0/g1_U_0 (.y ( f_out[4] ) , .b ( s1_start ) , .a ( \f_dout_master/genblk1[4].g0/n1 ));
  srdreg  \dout_master/genblk1[5].g0/g0_U (.ackout ( n1_N_3 ) , .f_q ( \f_dout_master/genblk1[5].g0/n1 ) , .t_q ( \t_dout_master/genblk1[5].g0/n1 ) , .f_d ( f_next_out[5] ) , .t_d ( t_next_out[5] ));
  and2  \dout_master/genblk1[5].g0/g1_U (.y ( t_out[5] ) , .b ( s1_start ) , .a ( \t_dout_master/genblk1[5].g0/n1 ));
  and2  \dout_master/genblk1_5_.g0/g1_U_0 (.y ( f_out[5] ) , .b ( s1_start ) , .a ( \f_dout_master/genblk1[5].g0/n1 ));
  srdreg  \dout_master/genblk1[6].g0/g0_U (.ackout ( n1_N_4 ) , .f_q ( \f_dout_master/genblk1[6].g0/n1 ) , .t_q ( \t_dout_master/genblk1[6].g0/n1 ) , .f_d ( f_next_out[6] ) , .t_d ( t_next_out[6] ));
  and2  \dout_master/genblk1[6].g0/g1_U (.y ( t_out[6] ) , .b ( s1_start ) , .a ( \t_dout_master/genblk1[6].g0/n1 ));
  and2  \dout_master/genblk1_6_.g0/g1_U_0 (.y ( f_out[6] ) , .b ( s1_start ) , .a ( \f_dout_master/genblk1[6].g0/n1 ));
  srdreg  \dout_master/genblk1[7].g0/g0_U (.ackout ( n1_N_5 ) , .f_q ( \f_dout_master/genblk1[7].g0/n1 ) , .t_q ( \t_dout_master/genblk1[7].g0/n1 ) , .f_d ( f_next_out[7] ) , .t_d ( t_next_out[7] ));
  and2  \dout_master/genblk1[7].g0/g1_U (.y ( t_out[7] ) , .b ( s1_start ) , .a ( \t_dout_master/genblk1[7].g0/n1 ));
  and2  \dout_master/genblk1_7_.g0/g1_U_0 (.y ( f_out[7] ) , .b ( s1_start ) , .a ( \f_dout_master/genblk1[7].g0/n1 ));
  srdreg  \dout_slave/genblk1[0].g0/g0_U (.ackout ( n1_N_6 ) , .f_q ( \f_dout_slave/genblk1[0].g0/n1 ) , .t_q ( \t_dout_slave/genblk1[0].g0/n1 ) , .f_d ( f_out[0] ) , .t_d ( t_out[0] ));
  and2  \dout_slave/genblk1[0].g0/g1_U (.y ( t_out_now[0] ) , .b ( s0 ) , .a ( \t_dout_slave/genblk1[0].g0/n1 ));
  and2  \dout_slave/genblk1_0_.g0/g1_U_0 (.y ( f_out_now[0] ) , .b ( s0 ) , .a ( \f_dout_slave/genblk1[0].g0/n1 ));
  srdreg  \dout_slave/genblk1[1].g0/g0_U (.ackout ( n1_N_7 ) , .f_q ( \f_dout_slave/genblk1[1].g0/n1 ) , .t_q ( \t_dout_slave/genblk1[1].g0/n1 ) , .f_d ( f_out[1] ) , .t_d ( t_out[1] ));
  and2  \dout_slave/genblk1[1].g0/g1_U (.y ( t_out_now[1] ) , .b ( s0 ) , .a ( \t_dout_slave/genblk1[1].g0/n1 ));
  and2  \dout_slave/genblk1_1_.g0/g1_U_0 (.y ( f_out_now[1] ) , .b ( s0 ) , .a ( \f_dout_slave/genblk1[1].g0/n1 ));
  srdreg  \dout_slave/genblk1[2].g0/g0_U (.ackout ( n1_N_8 ) , .f_q ( \f_dout_slave/genblk1[2].g0/n1 ) , .t_q ( \t_dout_slave/genblk1[2].g0/n1 ) , .f_d ( f_out[2] ) , .t_d ( t_out[2] ));
  and2  \dout_slave/genblk1[2].g0/g1_U (.y ( t_out_now[2] ) , .b ( s0 ) , .a ( \t_dout_slave/genblk1[2].g0/n1 ));
  and2  \dout_slave/genblk1_2_.g0/g1_U_0 (.y ( f_out_now[2] ) , .b ( s0 ) , .a ( \f_dout_slave/genblk1[2].g0/n1 ));
  srdreg  \dout_slave/genblk1[3].g0/g0_U (.ackout ( n1_N_9 ) , .f_q ( \f_dout_slave/genblk1[3].g0/n1 ) , .t_q ( \t_dout_slave/genblk1[3].g0/n1 ) , .f_d ( f_out[3] ) , .t_d ( t_out[3] ));
  and2  \dout_slave/genblk1[3].g0/g1_U (.y ( t_out_now[3] ) , .b ( s0 ) , .a ( \t_dout_slave/genblk1[3].g0/n1 ));
  and2  \dout_slave/genblk1_3_.g0/g1_U_0 (.y ( f_out_now[3] ) , .b ( s0 ) , .a ( \f_dout_slave/genblk1[3].g0/n1 ));
  srdreg  \dout_slave/genblk1[4].g0/g0_U (.ackout ( n1_N_10 ) , .f_q ( \f_dout_slave/genblk1[4].g0/n1 ) , .t_q ( \t_dout_slave/genblk1[4].g0/n1 ) , .f_d ( f_out[4] ) , .t_d ( t_out[4] ));
  and2  \dout_slave/genblk1[4].g0/g1_U (.y ( t_out_now[4] ) , .b ( s0 ) , .a ( \t_dout_slave/genblk1[4].g0/n1 ));
  and2  \dout_slave/genblk1_4_.g0/g1_U_0 (.y ( f_out_now[4] ) , .b ( s0 ) , .a ( \f_dout_slave/genblk1[4].g0/n1 ));
  srdreg  \dout_slave/genblk1[5].g0/g0_U (.ackout ( n1_N_11 ) , .f_q ( \f_dout_slave/genblk1[5].g0/n1 ) , .t_q ( \t_dout_slave/genblk1[5].g0/n1 ) , .f_d ( f_out[5] ) , .t_d ( t_out[5] ));
  and2  \dout_slave/genblk1[5].g0/g1_U (.y ( t_out_now[5] ) , .b ( s0 ) , .a ( \t_dout_slave/genblk1[5].g0/n1 ));
  and2  \dout_slave/genblk1_5_.g0/g1_U_0 (.y ( f_out_now[5] ) , .b ( s0 ) , .a ( \f_dout_slave/genblk1[5].g0/n1 ));
  srdreg  \dout_slave/genblk1[6].g0/g0_U (.ackout ( n1_N_12 ) , .f_q ( \f_dout_slave/genblk1[6].g0/n1 ) , .t_q ( \t_dout_slave/genblk1[6].g0/n1 ) , .f_d ( f_out[6] ) , .t_d ( t_out[6] ));
  and2  \dout_slave/genblk1[6].g0/g1_U (.y ( t_out_now[6] ) , .b ( s0 ) , .a ( \t_dout_slave/genblk1[6].g0/n1 ));
  and2  \dout_slave/genblk1_6_.g0/g1_U_0 (.y ( f_out_now[6] ) , .b ( s0 ) , .a ( \f_dout_slave/genblk1[6].g0/n1 ));
  srdreg  \dout_slave/genblk1[7].g0/g0_U (.ackout ( n1_N_13 ) , .f_q ( \f_dout_slave/genblk1[7].g0/n1 ) , .t_q ( \t_dout_slave/genblk1[7].g0/n1 ) , .f_d ( f_out[7] ) , .t_d ( t_out[7] ));
  and2  \dout_slave/genblk1[7].g0/g1_U (.y ( t_out_now[7] ) , .b ( s0 ) , .a ( \t_dout_slave/genblk1[7].g0/n1 ));
  and2  \dout_slave/genblk1_7_.g0/g1_U_0 (.y ( f_out_now[7] ) , .b ( s0 ) , .a ( \f_dout_slave/genblk1[7].g0/n1 ));
  srdreg  \dout_master/genblk1[0].g0/g0_U (.ackout ( n1_N_14 ) , .f_q ( \f_dout_master/genblk1[0].g0/n1 ) , .t_q ( \t_dout_master/genblk1[0].g0/n1 ) , .f_d ( f_next_out[0] ) , .t_d ( t_next_out[0] ));
  and2  \dout_master/genblk1[0].g0/g1_U (.y ( t_out[0] ) , .b ( s1_start ) , .a ( \t_dout_master/genblk1[0].g0/n1 ));
  and2  \dout_master/genblk1_0_.g0/g1_U_0 (.y ( f_out[0] ) , .b ( s1_start ) , .a ( \f_dout_master/genblk1[0].g0/n1 ));
  thand0  U28_U (.y ( f_n4 ) , .d ( f_clr ) , .c ( f_enable ) , .b ( t_clr ) , .a ( t_enable ));
  th22  U28_U_0 (.y ( t_n4 ) , .b ( f_clr ) , .a ( f_enable ));
  thand0  U27_U (.y ( f_n17 ) , .d ( t_n4 ) , .c ( t_out_now[0] ) , .b ( f_n4 ) , .a ( f_out_now[0] ));
  th22  U27_U_0 (.y ( t_n17 ) , .b ( t_n4 ) , .a ( t_out_now[0] ));
  thand0  U26_U (.y ( f_n3 ) , .d ( t_enable ) , .c ( f_clr ) , .b ( f_enable ) , .a ( t_clr ));
  th22  U26_U_0 (.y ( t_n3 ) , .b ( t_enable ) , .a ( f_clr ));
  thand0  U25_U (.y ( f_n18 ) , .d ( t_n3 ) , .c ( f_out_now[0] ) , .b ( f_n3 ) , .a ( t_out_now[0] ));
  th22  U25_U_0 (.y ( t_n18 ) , .b ( t_n3 ) , .a ( f_out_now[0] ));
  thand0  U24_U (.y ( t_next_out[0] ) , .d ( f_n18 ) , .c ( f_n17 ) , .b ( t_n18 ) , .a ( t_n17 ));
  th22  U24_U_0 (.y ( f_next_out[0] ) , .b ( f_n18 ) , .a ( f_n17 ));
  thand0  U23_U (.y ( f_n15 ) , .d ( t_n4 ) , .c ( t_out_now[1] ) , .b ( f_n4 ) , .a ( f_out_now[1] ));
  th22  U23_U_0 (.y ( t_n15 ) , .b ( t_n4 ) , .a ( t_out_now[1] ));
  thand0  U22_U (.y ( f_n16 ) , .d ( t_n3 ) , .c ( t_N6 ) , .b ( f_n3 ) , .a ( f_N6 ));
  th22  U22_U_0 (.y ( t_n16 ) , .b ( t_n3 ) , .a ( t_N6 ));
  thand0  U21_U (.y ( t_next_out[1] ) , .d ( f_n16 ) , .c ( f_n15 ) , .b ( t_n16 ) , .a ( t_n15 ));
  th22  U21_U_0 (.y ( f_next_out[1] ) , .b ( f_n16 ) , .a ( f_n15 ));
  thand0  U20_U (.y ( f_n13 ) , .d ( t_n4 ) , .c ( t_out_now[2] ) , .b ( f_n4 ) , .a ( f_out_now[2] ));
  th22  U20_U_0 (.y ( t_n13 ) , .b ( t_n4 ) , .a ( t_out_now[2] ));
  thand0  U19_U (.y ( f_n14 ) , .d ( t_n3 ) , .c ( t_N7 ) , .b ( f_n3 ) , .a ( f_N7 ));
  th22  U19_U_0 (.y ( t_n14 ) , .b ( t_n3 ) , .a ( t_N7 ));
  thand0  U18_U (.y ( t_next_out[2] ) , .d ( f_n14 ) , .c ( f_n13 ) , .b ( t_n14 ) , .a ( t_n13 ));
  th22  U18_U_0 (.y ( f_next_out[2] ) , .b ( f_n14 ) , .a ( f_n13 ));
  thand0  U17_U (.y ( f_n11 ) , .d ( t_n4 ) , .c ( t_out_now[3] ) , .b ( f_n4 ) , .a ( f_out_now[3] ));
  th22  U17_U_0 (.y ( t_n11 ) , .b ( t_n4 ) , .a ( t_out_now[3] ));
  thand0  U16_U (.y ( f_n12 ) , .d ( t_n3 ) , .c ( t_N8 ) , .b ( f_n3 ) , .a ( f_N8 ));
  th22  U16_U_0 (.y ( t_n12 ) , .b ( t_n3 ) , .a ( t_N8 ));
  thand0  U15_U (.y ( t_next_out[3] ) , .d ( f_n12 ) , .c ( f_n11 ) , .b ( t_n12 ) , .a ( t_n11 ));
  th22  U15_U_0 (.y ( f_next_out[3] ) , .b ( f_n12 ) , .a ( f_n11 ));
  thand0  U14_U (.y ( f_n9 ) , .d ( t_n4 ) , .c ( t_out_now[4] ) , .b ( f_n4 ) , .a ( f_out_now[4] ));
  th22  U14_U_0 (.y ( t_n9 ) , .b ( t_n4 ) , .a ( t_out_now[4] ));
  thand0  U13_U (.y ( f_n10 ) , .d ( t_n3 ) , .c ( t_N9 ) , .b ( f_n3 ) , .a ( f_N9 ));
  th22  U13_U_0 (.y ( t_n10 ) , .b ( t_n3 ) , .a ( t_N9 ));
  thand0  U12_U (.y ( t_next_out[4] ) , .d ( f_n10 ) , .c ( f_n9 ) , .b ( t_n10 ) , .a ( t_n9 ));
  th22  U12_U_0 (.y ( f_next_out[4] ) , .b ( f_n10 ) , .a ( f_n9 ));
  thand0  U11_U (.y ( f_n7 ) , .d ( t_n4 ) , .c ( t_out_now[5] ) , .b ( f_n4 ) , .a ( f_out_now[5] ));
  th22  U11_U_0 (.y ( t_n7 ) , .b ( t_n4 ) , .a ( t_out_now[5] ));
  thand0  U10_U (.y ( f_n8 ) , .d ( t_n3 ) , .c ( t_N10 ) , .b ( f_n3 ) , .a ( f_N10 ));
  th22  U10_U_0 (.y ( t_n8 ) , .b ( t_n3 ) , .a ( t_N10 ));
  thand0  U9_U (.y ( t_next_out[5] ) , .d ( f_n8 ) , .c ( f_n7 ) , .b ( t_n8 ) , .a ( t_n7 ));
  th22  U9_U_0 (.y ( f_next_out[5] ) , .b ( f_n8 ) , .a ( f_n7 ));
  thand0  U8_U (.y ( f_n5 ) , .d ( t_n4 ) , .c ( t_out_now[6] ) , .b ( f_n4 ) , .a ( f_out_now[6] ));
  th22  U8_U_0 (.y ( t_n5 ) , .b ( t_n4 ) , .a ( t_out_now[6] ));
  thand0  U7_U (.y ( f_n6 ) , .d ( t_n3 ) , .c ( t_N11 ) , .b ( f_n3 ) , .a ( f_N11 ));
  th22  U7_U_0 (.y ( t_n6 ) , .b ( t_n3 ) , .a ( t_N11 ));
  thand0  U6_U (.y ( t_next_out[6] ) , .d ( f_n6 ) , .c ( f_n5 ) , .b ( t_n6 ) , .a ( t_n5 ));
  th22  U6_U_0 (.y ( f_next_out[6] ) , .b ( f_n6 ) , .a ( f_n5 ));
  thand0  U5_U (.y ( f_n1 ) , .d ( t_n4 ) , .c ( t_out_now[7] ) , .b ( f_n4 ) , .a ( f_out_now[7] ));
  th22  U5_U_0 (.y ( t_n1 ) , .b ( t_n4 ) , .a ( t_out_now[7] ));
  thand0  U4_U (.y ( f_n2 ) , .d ( t_n3 ) , .c ( t_N12 ) , .b ( f_n3 ) , .a ( f_N12 ));
  th22  U4_U_0 (.y ( t_n2 ) , .b ( t_n3 ) , .a ( t_N12 ));
  thand0  U3_U (.y ( t_next_out[7] ) , .d ( f_n2 ) , .c ( f_n1 ) , .b ( t_n2 ) , .a ( t_n1 ));
  th22  U3_U_0 (.y ( f_next_out[7] ) , .b ( f_n2 ) , .a ( f_n1 ));
  nor2  g0_U (.y ( s0_start ) , .b ( ki_N_0 ) , .a ( en_b_N ));
  inv  g0_U_0 (.y ( en_b_N ) , .a ( reset ));
endmodule
