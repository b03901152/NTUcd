//Unsigned 32x32=64 booth multiplier


module xnor2 (y, a, b);
output y;
input a,b;

wire yn;
xor2 g0 (.y(yn),.a(a),.b(b));
inv g1 (.y(y),.a(yn));
endmodule

module and3 (y, a, b, c);
output y;
input a,b,c;

wire n1;
and2 g0 (.y(n1),.a(a),.b(b));
and2 g1 (.y(y),.a(n1),.b(c));
endmodule


module ha(s,co,a,b);
output s,co;
input a,b;

and2 g0 (.y(co),.a(a),.b(b));
xor2 g1 (.y(s),.a(a),.b(b));

endmodule


// xn = n2i+1, xc = x2i, xp = 
module booth_enc (xo,xo2,mo,xn,xc,xp);
output xo,xo2,mo;
input xn,xc,xp;

xor2 u0 (.y(xo),.a(xp), .b(xc));
inv  u1 (.y(xn_b),.a(xn));
inv  u2 (.y(xc_b),.a(xc));
inv  u3 (.y(xp_b),.a(xp));
and3 u4 (.y(n1),.a(xp), .b(xc),.c(xn_b));
and3 u5 (.y(n2),.a(xp_b), .b(xc_b),.c(xn));
or2 u6 (.y(xo2),.a(n1),.b(n2));

assign mo = xn;

endmodule


module booth_sel (p,y1,y0,x2,x,m);
output p;
input y1,y0,x2,x,m;

and2 g0 (.y(nb),.a(y1),.b(x));
and2 g1 (.y(na),.a(y0),.b(x2));
or2 g2 (.y(nc),.a(nb),.b(na));
inv g3(.y(n1),.a(nc));

xnor2 u1 (.y(p), .a(n1),.b(m));
endmodule



module mult32x32 (a,b,p);

input [31:0] a,b;
output [63:0] p;

wire [47:0] s_vec,c_vec;
wire [32:0] a_int,b_int;
wire co0_0;
wire co1_0;
wire co2_0;
wire co3_0;
wire co4_0;
wire co5_0;
wire co6_0;
wire co7_0;
wire co8_0;
wire co9_0;
wire co10_0;
wire co11_0;
wire co12_0;
wire co13_0;
wire co14_0;
wire co15_0;
wire co16_0;
assign sig0 = 0;
assign sig1 = 1;
assign a_int[31:0] = a;
assign b_int[31:0] = b;
assign a_int[32] = sig0;
assign b_int[32] = sig0;
//Booth Select: 0
  booth_enc u_benc_0 (.xo(xo_0),.xo2(xo2_0),.mo(mo_0),.xn(a_int[1]),.xc(a_int[0]),.xp(sig0));
  inv u_mo0_n (.y(mo0_n),.a(mo_0));
  assign sbit0 = mo_0;
  assign sbit0_n = mo0_n;
  booth_sel u_pp0_0 (.p(pp0_0),.y1(b_int[0]),.y0(sig0),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_1 (.p(pp0_1),.y1(b_int[1]),.y0(b_int[0]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_2 (.p(pp0_2),.y1(b_int[2]),.y0(b_int[1]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_3 (.p(pp0_3),.y1(b_int[3]),.y0(b_int[2]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_4 (.p(pp0_4),.y1(b_int[4]),.y0(b_int[3]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_5 (.p(pp0_5),.y1(b_int[5]),.y0(b_int[4]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_6 (.p(pp0_6),.y1(b_int[6]),.y0(b_int[5]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_7 (.p(pp0_7),.y1(b_int[7]),.y0(b_int[6]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_8 (.p(pp0_8),.y1(b_int[8]),.y0(b_int[7]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_9 (.p(pp0_9),.y1(b_int[9]),.y0(b_int[8]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_10 (.p(pp0_10),.y1(b_int[10]),.y0(b_int[9]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_11 (.p(pp0_11),.y1(b_int[11]),.y0(b_int[10]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_12 (.p(pp0_12),.y1(b_int[12]),.y0(b_int[11]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_13 (.p(pp0_13),.y1(b_int[13]),.y0(b_int[12]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_14 (.p(pp0_14),.y1(b_int[14]),.y0(b_int[13]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_15 (.p(pp0_15),.y1(b_int[15]),.y0(b_int[14]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_16 (.p(pp0_16),.y1(b_int[16]),.y0(b_int[15]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_17 (.p(pp0_17),.y1(b_int[17]),.y0(b_int[16]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_18 (.p(pp0_18),.y1(b_int[18]),.y0(b_int[17]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_19 (.p(pp0_19),.y1(b_int[19]),.y0(b_int[18]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_20 (.p(pp0_20),.y1(b_int[20]),.y0(b_int[19]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_21 (.p(pp0_21),.y1(b_int[21]),.y0(b_int[20]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_22 (.p(pp0_22),.y1(b_int[22]),.y0(b_int[21]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_23 (.p(pp0_23),.y1(b_int[23]),.y0(b_int[22]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_24 (.p(pp0_24),.y1(b_int[24]),.y0(b_int[23]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_25 (.p(pp0_25),.y1(b_int[25]),.y0(b_int[24]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_26 (.p(pp0_26),.y1(b_int[26]),.y0(b_int[25]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_27 (.p(pp0_27),.y1(b_int[27]),.y0(b_int[26]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_28 (.p(pp0_28),.y1(b_int[28]),.y0(b_int[27]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_29 (.p(pp0_29),.y1(b_int[29]),.y0(b_int[28]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_30 (.p(pp0_30),.y1(b_int[30]),.y0(b_int[29]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_31 (.p(pp0_31),.y1(b_int[31]),.y0(b_int[30]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  booth_sel u_pp0_32 (.p(pp0_32),.y1(b_int[32]),.y0(b_int[31]),.x(xo_0),.x2(xo2_0),.m(mo_0));
  assign pp0_33 = sbit0;
  assign pp0_34 = sbit0;
  assign pp0_35 = sbit0_n;
//Booth Select: 1
  booth_enc u_benc_1 (.xo(xo_1),.xo2(xo2_1),.mo(mo_1),.xn(a_int[3]),.xc(a_int[2]),.xp(a_int[1]));
  inv u_mo1_n (.y(mo1_n),.a(mo_1));
  assign sbit1 = mo_1;
  assign sbit1_n = mo1_n;
  assign pp1_0 = sbit0;
  assign pp1_1 = sig0;
  booth_sel u_pp1_2 (.p(pp1_2),.y1(b_int[0]),.y0(sig0),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_3 (.p(pp1_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_4 (.p(pp1_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_5 (.p(pp1_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_6 (.p(pp1_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_7 (.p(pp1_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_8 (.p(pp1_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_9 (.p(pp1_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_10 (.p(pp1_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_11 (.p(pp1_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_12 (.p(pp1_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_13 (.p(pp1_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_14 (.p(pp1_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_15 (.p(pp1_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_16 (.p(pp1_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_17 (.p(pp1_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_18 (.p(pp1_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_19 (.p(pp1_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_20 (.p(pp1_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_21 (.p(pp1_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_22 (.p(pp1_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_23 (.p(pp1_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_24 (.p(pp1_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_25 (.p(pp1_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_26 (.p(pp1_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_27 (.p(pp1_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_28 (.p(pp1_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_29 (.p(pp1_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_30 (.p(pp1_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_31 (.p(pp1_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_32 (.p(pp1_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_33 (.p(pp1_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  booth_sel u_pp1_34 (.p(pp1_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_1),.x2(xo2_1),.m(mo_1));
  assign pp1_35 = sbit1_n;
  assign pp1_36 = sig1;
//Booth Select: 2
  booth_enc u_benc_2 (.xo(xo_2),.xo2(xo2_2),.mo(mo_2),.xn(a_int[5]),.xc(a_int[4]),.xp(a_int[3]));
  inv u_mo2_n (.y(mo2_n),.a(mo_2));
  assign sbit2 = mo_2;
  assign sbit2_n = mo2_n;
  assign pp2_0 = sbit1;
  assign pp2_1 = sig0;
  booth_sel u_pp2_2 (.p(pp2_2),.y1(b_int[0]),.y0(sig0),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_3 (.p(pp2_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_4 (.p(pp2_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_5 (.p(pp2_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_6 (.p(pp2_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_7 (.p(pp2_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_8 (.p(pp2_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_9 (.p(pp2_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_10 (.p(pp2_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_11 (.p(pp2_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_12 (.p(pp2_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_13 (.p(pp2_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_14 (.p(pp2_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_15 (.p(pp2_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_16 (.p(pp2_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_17 (.p(pp2_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_18 (.p(pp2_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_19 (.p(pp2_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_20 (.p(pp2_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_21 (.p(pp2_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_22 (.p(pp2_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_23 (.p(pp2_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_24 (.p(pp2_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_25 (.p(pp2_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_26 (.p(pp2_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_27 (.p(pp2_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_28 (.p(pp2_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_29 (.p(pp2_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_30 (.p(pp2_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_31 (.p(pp2_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_32 (.p(pp2_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_33 (.p(pp2_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  booth_sel u_pp2_34 (.p(pp2_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_2),.x2(xo2_2),.m(mo_2));
  assign pp2_35 = sbit2_n;
  assign pp2_36 = sig1;
//Booth Select: 3
  booth_enc u_benc_3 (.xo(xo_3),.xo2(xo2_3),.mo(mo_3),.xn(a_int[7]),.xc(a_int[6]),.xp(a_int[5]));
  inv u_mo3_n (.y(mo3_n),.a(mo_3));
  assign sbit3 = mo_3;
  assign sbit3_n = mo3_n;
  assign pp3_0 = sbit2;
  assign pp3_1 = sig0;
  booth_sel u_pp3_2 (.p(pp3_2),.y1(b_int[0]),.y0(sig0),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_3 (.p(pp3_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_4 (.p(pp3_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_5 (.p(pp3_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_6 (.p(pp3_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_7 (.p(pp3_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_8 (.p(pp3_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_9 (.p(pp3_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_10 (.p(pp3_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_11 (.p(pp3_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_12 (.p(pp3_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_13 (.p(pp3_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_14 (.p(pp3_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_15 (.p(pp3_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_16 (.p(pp3_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_17 (.p(pp3_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_18 (.p(pp3_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_19 (.p(pp3_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_20 (.p(pp3_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_21 (.p(pp3_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_22 (.p(pp3_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_23 (.p(pp3_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_24 (.p(pp3_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_25 (.p(pp3_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_26 (.p(pp3_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_27 (.p(pp3_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_28 (.p(pp3_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_29 (.p(pp3_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_30 (.p(pp3_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_31 (.p(pp3_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_32 (.p(pp3_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_33 (.p(pp3_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  booth_sel u_pp3_34 (.p(pp3_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_3),.x2(xo2_3),.m(mo_3));
  assign pp3_35 = sbit3_n;
  assign pp3_36 = sig1;
//Booth Select: 4
  booth_enc u_benc_4 (.xo(xo_4),.xo2(xo2_4),.mo(mo_4),.xn(a_int[9]),.xc(a_int[8]),.xp(a_int[7]));
  inv u_mo4_n (.y(mo4_n),.a(mo_4));
  assign sbit4 = mo_4;
  assign sbit4_n = mo4_n;
  assign pp4_0 = sbit3;
  assign pp4_1 = sig0;
  booth_sel u_pp4_2 (.p(pp4_2),.y1(b_int[0]),.y0(sig0),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_3 (.p(pp4_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_4 (.p(pp4_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_5 (.p(pp4_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_6 (.p(pp4_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_7 (.p(pp4_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_8 (.p(pp4_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_9 (.p(pp4_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_10 (.p(pp4_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_11 (.p(pp4_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_12 (.p(pp4_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_13 (.p(pp4_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_14 (.p(pp4_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_15 (.p(pp4_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_16 (.p(pp4_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_17 (.p(pp4_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_18 (.p(pp4_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_19 (.p(pp4_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_20 (.p(pp4_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_21 (.p(pp4_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_22 (.p(pp4_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_23 (.p(pp4_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_24 (.p(pp4_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_25 (.p(pp4_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_26 (.p(pp4_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_27 (.p(pp4_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_28 (.p(pp4_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_29 (.p(pp4_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_30 (.p(pp4_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_31 (.p(pp4_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_32 (.p(pp4_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_33 (.p(pp4_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  booth_sel u_pp4_34 (.p(pp4_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_4),.x2(xo2_4),.m(mo_4));
  assign pp4_35 = sbit4_n;
  assign pp4_36 = sig1;
//Booth Select: 5
  booth_enc u_benc_5 (.xo(xo_5),.xo2(xo2_5),.mo(mo_5),.xn(a_int[11]),.xc(a_int[10]),.xp(a_int[9]));
  inv u_mo5_n (.y(mo5_n),.a(mo_5));
  assign sbit5 = mo_5;
  assign sbit5_n = mo5_n;
  assign pp5_0 = sbit4;
  assign pp5_1 = sig0;
  booth_sel u_pp5_2 (.p(pp5_2),.y1(b_int[0]),.y0(sig0),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_3 (.p(pp5_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_4 (.p(pp5_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_5 (.p(pp5_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_6 (.p(pp5_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_7 (.p(pp5_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_8 (.p(pp5_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_9 (.p(pp5_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_10 (.p(pp5_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_11 (.p(pp5_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_12 (.p(pp5_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_13 (.p(pp5_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_14 (.p(pp5_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_15 (.p(pp5_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_16 (.p(pp5_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_17 (.p(pp5_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_18 (.p(pp5_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_19 (.p(pp5_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_20 (.p(pp5_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_21 (.p(pp5_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_22 (.p(pp5_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_23 (.p(pp5_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_24 (.p(pp5_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_25 (.p(pp5_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_26 (.p(pp5_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_27 (.p(pp5_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_28 (.p(pp5_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_29 (.p(pp5_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_30 (.p(pp5_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_31 (.p(pp5_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_32 (.p(pp5_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_33 (.p(pp5_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  booth_sel u_pp5_34 (.p(pp5_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_5),.x2(xo2_5),.m(mo_5));
  assign pp5_35 = sbit5_n;
  assign pp5_36 = sig1;
//Booth Select: 6
  booth_enc u_benc_6 (.xo(xo_6),.xo2(xo2_6),.mo(mo_6),.xn(a_int[13]),.xc(a_int[12]),.xp(a_int[11]));
  inv u_mo6_n (.y(mo6_n),.a(mo_6));
  assign sbit6 = mo_6;
  assign sbit6_n = mo6_n;
  assign pp6_0 = sbit5;
  assign pp6_1 = sig0;
  booth_sel u_pp6_2 (.p(pp6_2),.y1(b_int[0]),.y0(sig0),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_3 (.p(pp6_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_4 (.p(pp6_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_5 (.p(pp6_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_6 (.p(pp6_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_7 (.p(pp6_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_8 (.p(pp6_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_9 (.p(pp6_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_10 (.p(pp6_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_11 (.p(pp6_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_12 (.p(pp6_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_13 (.p(pp6_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_14 (.p(pp6_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_15 (.p(pp6_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_16 (.p(pp6_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_17 (.p(pp6_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_18 (.p(pp6_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_19 (.p(pp6_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_20 (.p(pp6_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_21 (.p(pp6_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_22 (.p(pp6_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_23 (.p(pp6_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_24 (.p(pp6_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_25 (.p(pp6_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_26 (.p(pp6_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_27 (.p(pp6_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_28 (.p(pp6_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_29 (.p(pp6_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_30 (.p(pp6_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_31 (.p(pp6_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_32 (.p(pp6_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_33 (.p(pp6_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  booth_sel u_pp6_34 (.p(pp6_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_6),.x2(xo2_6),.m(mo_6));
  assign pp6_35 = sbit6_n;
  assign pp6_36 = sig1;
//Booth Select: 7
  booth_enc u_benc_7 (.xo(xo_7),.xo2(xo2_7),.mo(mo_7),.xn(a_int[15]),.xc(a_int[14]),.xp(a_int[13]));
  inv u_mo7_n (.y(mo7_n),.a(mo_7));
  assign sbit7 = mo_7;
  assign sbit7_n = mo7_n;
  assign pp7_0 = sbit6;
  assign pp7_1 = sig0;
  booth_sel u_pp7_2 (.p(pp7_2),.y1(b_int[0]),.y0(sig0),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_3 (.p(pp7_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_4 (.p(pp7_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_5 (.p(pp7_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_6 (.p(pp7_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_7 (.p(pp7_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_8 (.p(pp7_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_9 (.p(pp7_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_10 (.p(pp7_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_11 (.p(pp7_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_12 (.p(pp7_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_13 (.p(pp7_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_14 (.p(pp7_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_15 (.p(pp7_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_16 (.p(pp7_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_17 (.p(pp7_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_18 (.p(pp7_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_19 (.p(pp7_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_20 (.p(pp7_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_21 (.p(pp7_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_22 (.p(pp7_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_23 (.p(pp7_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_24 (.p(pp7_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_25 (.p(pp7_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_26 (.p(pp7_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_27 (.p(pp7_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_28 (.p(pp7_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_29 (.p(pp7_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_30 (.p(pp7_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_31 (.p(pp7_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_32 (.p(pp7_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_33 (.p(pp7_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  booth_sel u_pp7_34 (.p(pp7_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_7),.x2(xo2_7),.m(mo_7));
  assign pp7_35 = sbit7_n;
  assign pp7_36 = sig1;
//Booth Select: 8
  booth_enc u_benc_8 (.xo(xo_8),.xo2(xo2_8),.mo(mo_8),.xn(a_int[17]),.xc(a_int[16]),.xp(a_int[15]));
  inv u_mo8_n (.y(mo8_n),.a(mo_8));
  assign sbit8 = mo_8;
  assign sbit8_n = mo8_n;
  assign pp8_0 = sbit7;
  assign pp8_1 = sig0;
  booth_sel u_pp8_2 (.p(pp8_2),.y1(b_int[0]),.y0(sig0),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_3 (.p(pp8_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_4 (.p(pp8_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_5 (.p(pp8_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_6 (.p(pp8_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_7 (.p(pp8_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_8 (.p(pp8_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_9 (.p(pp8_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_10 (.p(pp8_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_11 (.p(pp8_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_12 (.p(pp8_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_13 (.p(pp8_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_14 (.p(pp8_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_15 (.p(pp8_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_16 (.p(pp8_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_17 (.p(pp8_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_18 (.p(pp8_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_19 (.p(pp8_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_20 (.p(pp8_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_21 (.p(pp8_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_22 (.p(pp8_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_23 (.p(pp8_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_24 (.p(pp8_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_25 (.p(pp8_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_26 (.p(pp8_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_27 (.p(pp8_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_28 (.p(pp8_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_29 (.p(pp8_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_30 (.p(pp8_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_31 (.p(pp8_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_32 (.p(pp8_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_33 (.p(pp8_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  booth_sel u_pp8_34 (.p(pp8_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_8),.x2(xo2_8),.m(mo_8));
  assign pp8_35 = sbit8_n;
  assign pp8_36 = sig1;
//Booth Select: 9
  booth_enc u_benc_9 (.xo(xo_9),.xo2(xo2_9),.mo(mo_9),.xn(a_int[19]),.xc(a_int[18]),.xp(a_int[17]));
  inv u_mo9_n (.y(mo9_n),.a(mo_9));
  assign sbit9 = mo_9;
  assign sbit9_n = mo9_n;
  assign pp9_0 = sbit8;
  assign pp9_1 = sig0;
  booth_sel u_pp9_2 (.p(pp9_2),.y1(b_int[0]),.y0(sig0),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_3 (.p(pp9_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_4 (.p(pp9_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_5 (.p(pp9_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_6 (.p(pp9_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_7 (.p(pp9_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_8 (.p(pp9_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_9 (.p(pp9_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_10 (.p(pp9_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_11 (.p(pp9_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_12 (.p(pp9_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_13 (.p(pp9_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_14 (.p(pp9_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_15 (.p(pp9_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_16 (.p(pp9_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_17 (.p(pp9_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_18 (.p(pp9_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_19 (.p(pp9_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_20 (.p(pp9_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_21 (.p(pp9_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_22 (.p(pp9_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_23 (.p(pp9_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_24 (.p(pp9_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_25 (.p(pp9_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_26 (.p(pp9_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_27 (.p(pp9_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_28 (.p(pp9_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_29 (.p(pp9_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_30 (.p(pp9_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_31 (.p(pp9_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_32 (.p(pp9_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_33 (.p(pp9_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  booth_sel u_pp9_34 (.p(pp9_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_9),.x2(xo2_9),.m(mo_9));
  assign pp9_35 = sbit9_n;
  assign pp9_36 = sig1;
//Booth Select: 10
  booth_enc u_benc_10 (.xo(xo_10),.xo2(xo2_10),.mo(mo_10),.xn(a_int[21]),.xc(a_int[20]),.xp(a_int[19]));
  inv u_mo10_n (.y(mo10_n),.a(mo_10));
  assign sbit10 = mo_10;
  assign sbit10_n = mo10_n;
  assign pp10_0 = sbit9;
  assign pp10_1 = sig0;
  booth_sel u_pp10_2 (.p(pp10_2),.y1(b_int[0]),.y0(sig0),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_3 (.p(pp10_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_4 (.p(pp10_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_5 (.p(pp10_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_6 (.p(pp10_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_7 (.p(pp10_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_8 (.p(pp10_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_9 (.p(pp10_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_10 (.p(pp10_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_11 (.p(pp10_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_12 (.p(pp10_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_13 (.p(pp10_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_14 (.p(pp10_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_15 (.p(pp10_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_16 (.p(pp10_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_17 (.p(pp10_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_18 (.p(pp10_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_19 (.p(pp10_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_20 (.p(pp10_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_21 (.p(pp10_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_22 (.p(pp10_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_23 (.p(pp10_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_24 (.p(pp10_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_25 (.p(pp10_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_26 (.p(pp10_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_27 (.p(pp10_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_28 (.p(pp10_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_29 (.p(pp10_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_30 (.p(pp10_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_31 (.p(pp10_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_32 (.p(pp10_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_33 (.p(pp10_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  booth_sel u_pp10_34 (.p(pp10_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_10),.x2(xo2_10),.m(mo_10));
  assign pp10_35 = sbit10_n;
  assign pp10_36 = sig1;
//Booth Select: 11
  booth_enc u_benc_11 (.xo(xo_11),.xo2(xo2_11),.mo(mo_11),.xn(a_int[23]),.xc(a_int[22]),.xp(a_int[21]));
  inv u_mo11_n (.y(mo11_n),.a(mo_11));
  assign sbit11 = mo_11;
  assign sbit11_n = mo11_n;
  assign pp11_0 = sbit10;
  assign pp11_1 = sig0;
  booth_sel u_pp11_2 (.p(pp11_2),.y1(b_int[0]),.y0(sig0),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_3 (.p(pp11_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_4 (.p(pp11_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_5 (.p(pp11_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_6 (.p(pp11_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_7 (.p(pp11_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_8 (.p(pp11_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_9 (.p(pp11_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_10 (.p(pp11_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_11 (.p(pp11_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_12 (.p(pp11_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_13 (.p(pp11_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_14 (.p(pp11_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_15 (.p(pp11_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_16 (.p(pp11_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_17 (.p(pp11_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_18 (.p(pp11_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_19 (.p(pp11_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_20 (.p(pp11_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_21 (.p(pp11_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_22 (.p(pp11_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_23 (.p(pp11_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_24 (.p(pp11_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_25 (.p(pp11_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_26 (.p(pp11_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_27 (.p(pp11_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_28 (.p(pp11_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_29 (.p(pp11_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_30 (.p(pp11_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_31 (.p(pp11_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_32 (.p(pp11_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_33 (.p(pp11_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  booth_sel u_pp11_34 (.p(pp11_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_11),.x2(xo2_11),.m(mo_11));
  assign pp11_35 = sbit11_n;
  assign pp11_36 = sig1;
//Booth Select: 12
  booth_enc u_benc_12 (.xo(xo_12),.xo2(xo2_12),.mo(mo_12),.xn(a_int[25]),.xc(a_int[24]),.xp(a_int[23]));
  inv u_mo12_n (.y(mo12_n),.a(mo_12));
  assign sbit12 = mo_12;
  assign sbit12_n = mo12_n;
  assign pp12_0 = sbit11;
  assign pp12_1 = sig0;
  booth_sel u_pp12_2 (.p(pp12_2),.y1(b_int[0]),.y0(sig0),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_3 (.p(pp12_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_4 (.p(pp12_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_5 (.p(pp12_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_6 (.p(pp12_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_7 (.p(pp12_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_8 (.p(pp12_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_9 (.p(pp12_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_10 (.p(pp12_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_11 (.p(pp12_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_12 (.p(pp12_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_13 (.p(pp12_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_14 (.p(pp12_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_15 (.p(pp12_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_16 (.p(pp12_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_17 (.p(pp12_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_18 (.p(pp12_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_19 (.p(pp12_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_20 (.p(pp12_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_21 (.p(pp12_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_22 (.p(pp12_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_23 (.p(pp12_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_24 (.p(pp12_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_25 (.p(pp12_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_26 (.p(pp12_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_27 (.p(pp12_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_28 (.p(pp12_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_29 (.p(pp12_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_30 (.p(pp12_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_31 (.p(pp12_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_32 (.p(pp12_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_33 (.p(pp12_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  booth_sel u_pp12_34 (.p(pp12_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_12),.x2(xo2_12),.m(mo_12));
  assign pp12_35 = sbit12_n;
  assign pp12_36 = sig1;
//Booth Select: 13
  booth_enc u_benc_13 (.xo(xo_13),.xo2(xo2_13),.mo(mo_13),.xn(a_int[27]),.xc(a_int[26]),.xp(a_int[25]));
  inv u_mo13_n (.y(mo13_n),.a(mo_13));
  assign sbit13 = mo_13;
  assign sbit13_n = mo13_n;
  assign pp13_0 = sbit12;
  assign pp13_1 = sig0;
  booth_sel u_pp13_2 (.p(pp13_2),.y1(b_int[0]),.y0(sig0),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_3 (.p(pp13_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_4 (.p(pp13_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_5 (.p(pp13_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_6 (.p(pp13_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_7 (.p(pp13_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_8 (.p(pp13_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_9 (.p(pp13_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_10 (.p(pp13_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_11 (.p(pp13_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_12 (.p(pp13_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_13 (.p(pp13_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_14 (.p(pp13_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_15 (.p(pp13_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_16 (.p(pp13_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_17 (.p(pp13_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_18 (.p(pp13_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_19 (.p(pp13_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_20 (.p(pp13_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_21 (.p(pp13_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_22 (.p(pp13_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_23 (.p(pp13_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_24 (.p(pp13_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_25 (.p(pp13_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_26 (.p(pp13_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_27 (.p(pp13_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_28 (.p(pp13_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_29 (.p(pp13_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_30 (.p(pp13_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_31 (.p(pp13_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_32 (.p(pp13_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_33 (.p(pp13_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  booth_sel u_pp13_34 (.p(pp13_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_13),.x2(xo2_13),.m(mo_13));
  assign pp13_35 = sbit13_n;
  assign pp13_36 = sig1;
//Booth Select: 14
  booth_enc u_benc_14 (.xo(xo_14),.xo2(xo2_14),.mo(mo_14),.xn(a_int[29]),.xc(a_int[28]),.xp(a_int[27]));
  inv u_mo14_n (.y(mo14_n),.a(mo_14));
  assign sbit14 = mo_14;
  assign sbit14_n = mo14_n;
  assign pp14_0 = sbit13;
  assign pp14_1 = sig0;
  booth_sel u_pp14_2 (.p(pp14_2),.y1(b_int[0]),.y0(sig0),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_3 (.p(pp14_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_4 (.p(pp14_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_5 (.p(pp14_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_6 (.p(pp14_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_7 (.p(pp14_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_8 (.p(pp14_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_9 (.p(pp14_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_10 (.p(pp14_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_11 (.p(pp14_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_12 (.p(pp14_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_13 (.p(pp14_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_14 (.p(pp14_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_15 (.p(pp14_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_16 (.p(pp14_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_17 (.p(pp14_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_18 (.p(pp14_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_19 (.p(pp14_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_20 (.p(pp14_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_21 (.p(pp14_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_22 (.p(pp14_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_23 (.p(pp14_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_24 (.p(pp14_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_25 (.p(pp14_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_26 (.p(pp14_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_27 (.p(pp14_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_28 (.p(pp14_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_29 (.p(pp14_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_30 (.p(pp14_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_31 (.p(pp14_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_32 (.p(pp14_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_33 (.p(pp14_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  booth_sel u_pp14_34 (.p(pp14_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_14),.x2(xo2_14),.m(mo_14));
  assign pp14_35 = sbit14_n;
  assign pp14_36 = sig1;
//Booth Select: 15
  booth_enc u_benc_15 (.xo(xo_15),.xo2(xo2_15),.mo(mo_15),.xn(a_int[31]),.xc(a_int[30]),.xp(a_int[29]));
  inv u_mo15_n (.y(mo15_n),.a(mo_15));
  assign sbit15 = mo_15;
  assign sbit15_n = mo15_n;
  assign pp15_0 = sbit14;
  assign pp15_1 = sig0;
  booth_sel u_pp15_2 (.p(pp15_2),.y1(b_int[0]),.y0(sig0),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_3 (.p(pp15_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_4 (.p(pp15_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_5 (.p(pp15_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_6 (.p(pp15_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_7 (.p(pp15_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_8 (.p(pp15_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_9 (.p(pp15_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_10 (.p(pp15_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_11 (.p(pp15_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_12 (.p(pp15_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_13 (.p(pp15_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_14 (.p(pp15_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_15 (.p(pp15_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_16 (.p(pp15_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_17 (.p(pp15_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_18 (.p(pp15_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_19 (.p(pp15_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_20 (.p(pp15_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_21 (.p(pp15_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_22 (.p(pp15_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_23 (.p(pp15_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_24 (.p(pp15_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_25 (.p(pp15_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_26 (.p(pp15_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_27 (.p(pp15_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_28 (.p(pp15_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_29 (.p(pp15_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_30 (.p(pp15_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_31 (.p(pp15_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_32 (.p(pp15_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_33 (.p(pp15_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  booth_sel u_pp15_34 (.p(pp15_34),.y1(b_int[32]),.y0(b_int[31]),.x(xo_15),.x2(xo2_15),.m(mo_15));
  assign pp15_35 = sbit15_n;
//Booth Select: 16
  booth_enc u_benc_16 (.xo(xo_16),.xo2(xo2_16),.mo(mo_16),.xn(sig0),.xc(sig0),.xp(a_int[31]));
  assign pp16_0 = sbit15;
  assign pp16_1 = sig0;
  booth_sel u_pp16_2 (.p(pp16_2),.y1(b_int[0]),.y0(sig0),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_3 (.p(pp16_3),.y1(b_int[1]),.y0(b_int[0]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_4 (.p(pp16_4),.y1(b_int[2]),.y0(b_int[1]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_5 (.p(pp16_5),.y1(b_int[3]),.y0(b_int[2]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_6 (.p(pp16_6),.y1(b_int[4]),.y0(b_int[3]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_7 (.p(pp16_7),.y1(b_int[5]),.y0(b_int[4]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_8 (.p(pp16_8),.y1(b_int[6]),.y0(b_int[5]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_9 (.p(pp16_9),.y1(b_int[7]),.y0(b_int[6]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_10 (.p(pp16_10),.y1(b_int[8]),.y0(b_int[7]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_11 (.p(pp16_11),.y1(b_int[9]),.y0(b_int[8]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_12 (.p(pp16_12),.y1(b_int[10]),.y0(b_int[9]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_13 (.p(pp16_13),.y1(b_int[11]),.y0(b_int[10]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_14 (.p(pp16_14),.y1(b_int[12]),.y0(b_int[11]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_15 (.p(pp16_15),.y1(b_int[13]),.y0(b_int[12]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_16 (.p(pp16_16),.y1(b_int[14]),.y0(b_int[13]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_17 (.p(pp16_17),.y1(b_int[15]),.y0(b_int[14]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_18 (.p(pp16_18),.y1(b_int[16]),.y0(b_int[15]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_19 (.p(pp16_19),.y1(b_int[17]),.y0(b_int[16]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_20 (.p(pp16_20),.y1(b_int[18]),.y0(b_int[17]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_21 (.p(pp16_21),.y1(b_int[19]),.y0(b_int[18]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_22 (.p(pp16_22),.y1(b_int[20]),.y0(b_int[19]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_23 (.p(pp16_23),.y1(b_int[21]),.y0(b_int[20]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_24 (.p(pp16_24),.y1(b_int[22]),.y0(b_int[21]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_25 (.p(pp16_25),.y1(b_int[23]),.y0(b_int[22]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_26 (.p(pp16_26),.y1(b_int[24]),.y0(b_int[23]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_27 (.p(pp16_27),.y1(b_int[25]),.y0(b_int[24]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_28 (.p(pp16_28),.y1(b_int[26]),.y0(b_int[25]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_29 (.p(pp16_29),.y1(b_int[27]),.y0(b_int[26]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_30 (.p(pp16_30),.y1(b_int[28]),.y0(b_int[27]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_31 (.p(pp16_31),.y1(b_int[29]),.y0(b_int[28]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_32 (.p(pp16_32),.y1(b_int[30]),.y0(b_int[29]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  booth_sel u_pp16_33 (.p(pp16_33),.y1(b_int[31]),.y0(b_int[30]),.x(xo_16),.x2(xo2_16),.m(mo_16));
  //CSA Array 
  //CSA Row 0 
  ha u_csa0_0 (.s(sum0_0),.co(co0_0),.a(pp1_0),.b(pp0_0));
  ha u_csa0_1 (.s(sum0_1),.co(co0_1),.a(pp1_1),.b(pp0_1));
  ha u_csa0_2 (.s(sum0_2),.co(co0_2),.a(pp1_2),.b(pp0_2));
  ha u_csa0_3 (.s(sum0_3),.co(co0_3),.a(pp1_3),.b(pp0_3));
  ha u_csa0_4 (.s(sum0_4),.co(co0_4),.a(pp1_4),.b(pp0_4));
  ha u_csa0_5 (.s(sum0_5),.co(co0_5),.a(pp1_5),.b(pp0_5));
  ha u_csa0_6 (.s(sum0_6),.co(co0_6),.a(pp1_6),.b(pp0_6));
  ha u_csa0_7 (.s(sum0_7),.co(co0_7),.a(pp1_7),.b(pp0_7));
  ha u_csa0_8 (.s(sum0_8),.co(co0_8),.a(pp1_8),.b(pp0_8));
  ha u_csa0_9 (.s(sum0_9),.co(co0_9),.a(pp1_9),.b(pp0_9));
  ha u_csa0_10 (.s(sum0_10),.co(co0_10),.a(pp1_10),.b(pp0_10));
  ha u_csa0_11 (.s(sum0_11),.co(co0_11),.a(pp1_11),.b(pp0_11));
  ha u_csa0_12 (.s(sum0_12),.co(co0_12),.a(pp1_12),.b(pp0_12));
  ha u_csa0_13 (.s(sum0_13),.co(co0_13),.a(pp1_13),.b(pp0_13));
  ha u_csa0_14 (.s(sum0_14),.co(co0_14),.a(pp1_14),.b(pp0_14));
  ha u_csa0_15 (.s(sum0_15),.co(co0_15),.a(pp1_15),.b(pp0_15));
  ha u_csa0_16 (.s(sum0_16),.co(co0_16),.a(pp1_16),.b(pp0_16));
  ha u_csa0_17 (.s(sum0_17),.co(co0_17),.a(pp1_17),.b(pp0_17));
  ha u_csa0_18 (.s(sum0_18),.co(co0_18),.a(pp1_18),.b(pp0_18));
  ha u_csa0_19 (.s(sum0_19),.co(co0_19),.a(pp1_19),.b(pp0_19));
  ha u_csa0_20 (.s(sum0_20),.co(co0_20),.a(pp1_20),.b(pp0_20));
  ha u_csa0_21 (.s(sum0_21),.co(co0_21),.a(pp1_21),.b(pp0_21));
  ha u_csa0_22 (.s(sum0_22),.co(co0_22),.a(pp1_22),.b(pp0_22));
  ha u_csa0_23 (.s(sum0_23),.co(co0_23),.a(pp1_23),.b(pp0_23));
  ha u_csa0_24 (.s(sum0_24),.co(co0_24),.a(pp1_24),.b(pp0_24));
  ha u_csa0_25 (.s(sum0_25),.co(co0_25),.a(pp1_25),.b(pp0_25));
  ha u_csa0_26 (.s(sum0_26),.co(co0_26),.a(pp1_26),.b(pp0_26));
  ha u_csa0_27 (.s(sum0_27),.co(co0_27),.a(pp1_27),.b(pp0_27));
  ha u_csa0_28 (.s(sum0_28),.co(co0_28),.a(pp1_28),.b(pp0_28));
  ha u_csa0_29 (.s(sum0_29),.co(co0_29),.a(pp1_29),.b(pp0_29));
  ha u_csa0_30 (.s(sum0_30),.co(co0_30),.a(pp1_30),.b(pp0_30));
  ha u_csa0_31 (.s(sum0_31),.co(co0_31),.a(pp1_31),.b(pp0_31));
  ha u_csa0_32 (.s(sum0_32),.co(co0_32),.a(pp1_32),.b(pp0_32));
  ha u_csa0_33 (.s(sum0_33),.co(co0_33),.a(pp1_33),.b(pp0_33));
  ha u_csa0_34 (.s(sum0_34),.co(co0_34),.a(pp1_34),.b(pp0_34));
  ha u_csa0_35 (.s(sum0_35),.co(co0_35),.a(pp1_35),.b(pp0_35));
  assign sum0_36=pp1_36;
  //CSA Row 1 
  ha u_csa1_0 (.s(sum1_0),.co(co1_0),.a(sum0_1),.b(co0_0));
  fa u_csa1_1 (.s(sum1_1),.co(co1_1),.a(pp2_0),.b(sum0_2),.ci(co0_1));
  fa u_csa1_2 (.s(sum1_2),.co(co1_2),.a(pp2_1),.b(sum0_3),.ci(co0_2));
  fa u_csa1_3 (.s(sum1_3),.co(co1_3),.a(pp2_2),.b(sum0_4),.ci(co0_3));
  fa u_csa1_4 (.s(sum1_4),.co(co1_4),.a(pp2_3),.b(sum0_5),.ci(co0_4));
  fa u_csa1_5 (.s(sum1_5),.co(co1_5),.a(pp2_4),.b(sum0_6),.ci(co0_5));
  fa u_csa1_6 (.s(sum1_6),.co(co1_6),.a(pp2_5),.b(sum0_7),.ci(co0_6));
  fa u_csa1_7 (.s(sum1_7),.co(co1_7),.a(pp2_6),.b(sum0_8),.ci(co0_7));
  fa u_csa1_8 (.s(sum1_8),.co(co1_8),.a(pp2_7),.b(sum0_9),.ci(co0_8));
  fa u_csa1_9 (.s(sum1_9),.co(co1_9),.a(pp2_8),.b(sum0_10),.ci(co0_9));
  fa u_csa1_10 (.s(sum1_10),.co(co1_10),.a(pp2_9),.b(sum0_11),.ci(co0_10));
  fa u_csa1_11 (.s(sum1_11),.co(co1_11),.a(pp2_10),.b(sum0_12),.ci(co0_11));
  fa u_csa1_12 (.s(sum1_12),.co(co1_12),.a(pp2_11),.b(sum0_13),.ci(co0_12));
  fa u_csa1_13 (.s(sum1_13),.co(co1_13),.a(pp2_12),.b(sum0_14),.ci(co0_13));
  fa u_csa1_14 (.s(sum1_14),.co(co1_14),.a(pp2_13),.b(sum0_15),.ci(co0_14));
  fa u_csa1_15 (.s(sum1_15),.co(co1_15),.a(pp2_14),.b(sum0_16),.ci(co0_15));
  fa u_csa1_16 (.s(sum1_16),.co(co1_16),.a(pp2_15),.b(sum0_17),.ci(co0_16));
  fa u_csa1_17 (.s(sum1_17),.co(co1_17),.a(pp2_16),.b(sum0_18),.ci(co0_17));
  fa u_csa1_18 (.s(sum1_18),.co(co1_18),.a(pp2_17),.b(sum0_19),.ci(co0_18));
  fa u_csa1_19 (.s(sum1_19),.co(co1_19),.a(pp2_18),.b(sum0_20),.ci(co0_19));
  fa u_csa1_20 (.s(sum1_20),.co(co1_20),.a(pp2_19),.b(sum0_21),.ci(co0_20));
  fa u_csa1_21 (.s(sum1_21),.co(co1_21),.a(pp2_20),.b(sum0_22),.ci(co0_21));
  fa u_csa1_22 (.s(sum1_22),.co(co1_22),.a(pp2_21),.b(sum0_23),.ci(co0_22));
  fa u_csa1_23 (.s(sum1_23),.co(co1_23),.a(pp2_22),.b(sum0_24),.ci(co0_23));
  fa u_csa1_24 (.s(sum1_24),.co(co1_24),.a(pp2_23),.b(sum0_25),.ci(co0_24));
  fa u_csa1_25 (.s(sum1_25),.co(co1_25),.a(pp2_24),.b(sum0_26),.ci(co0_25));
  fa u_csa1_26 (.s(sum1_26),.co(co1_26),.a(pp2_25),.b(sum0_27),.ci(co0_26));
  fa u_csa1_27 (.s(sum1_27),.co(co1_27),.a(pp2_26),.b(sum0_28),.ci(co0_27));
  fa u_csa1_28 (.s(sum1_28),.co(co1_28),.a(pp2_27),.b(sum0_29),.ci(co0_28));
  fa u_csa1_29 (.s(sum1_29),.co(co1_29),.a(pp2_28),.b(sum0_30),.ci(co0_29));
  fa u_csa1_30 (.s(sum1_30),.co(co1_30),.a(pp2_29),.b(sum0_31),.ci(co0_30));
  fa u_csa1_31 (.s(sum1_31),.co(co1_31),.a(pp2_30),.b(sum0_32),.ci(co0_31));
  fa u_csa1_32 (.s(sum1_32),.co(co1_32),.a(pp2_31),.b(sum0_33),.ci(co0_32));
  fa u_csa1_33 (.s(sum1_33),.co(co1_33),.a(pp2_32),.b(sum0_34),.ci(co0_33));
  fa u_csa1_34 (.s(sum1_34),.co(co1_34),.a(pp2_33),.b(sum0_35),.ci(co0_34));
  fa u_csa1_35 (.s(sum1_35),.co(co1_35),.a(pp2_34),.b(sum0_36),.ci(co0_35));
  assign sum1_36=pp2_35;
  assign co1_36=sig0;
  assign sum1_37=pp2_36;
  //CSA Row 2 
  ha u_csa2_0 (.s(sum2_0),.co(co2_0),.a(sum1_1),.b(co1_0));
  ha u_csa2_1 (.s(sum2_1),.co(co2_1),.a(sum1_2),.b(co1_1));
  fa u_csa2_2 (.s(sum2_2),.co(co2_2),.a(pp3_0),.b(sum1_3),.ci(co1_2));
  fa u_csa2_3 (.s(sum2_3),.co(co2_3),.a(pp3_1),.b(sum1_4),.ci(co1_3));
  fa u_csa2_4 (.s(sum2_4),.co(co2_4),.a(pp3_2),.b(sum1_5),.ci(co1_4));
  fa u_csa2_5 (.s(sum2_5),.co(co2_5),.a(pp3_3),.b(sum1_6),.ci(co1_5));
  fa u_csa2_6 (.s(sum2_6),.co(co2_6),.a(pp3_4),.b(sum1_7),.ci(co1_6));
  fa u_csa2_7 (.s(sum2_7),.co(co2_7),.a(pp3_5),.b(sum1_8),.ci(co1_7));
  fa u_csa2_8 (.s(sum2_8),.co(co2_8),.a(pp3_6),.b(sum1_9),.ci(co1_8));
  fa u_csa2_9 (.s(sum2_9),.co(co2_9),.a(pp3_7),.b(sum1_10),.ci(co1_9));
  fa u_csa2_10 (.s(sum2_10),.co(co2_10),.a(pp3_8),.b(sum1_11),.ci(co1_10));
  fa u_csa2_11 (.s(sum2_11),.co(co2_11),.a(pp3_9),.b(sum1_12),.ci(co1_11));
  fa u_csa2_12 (.s(sum2_12),.co(co2_12),.a(pp3_10),.b(sum1_13),.ci(co1_12));
  fa u_csa2_13 (.s(sum2_13),.co(co2_13),.a(pp3_11),.b(sum1_14),.ci(co1_13));
  fa u_csa2_14 (.s(sum2_14),.co(co2_14),.a(pp3_12),.b(sum1_15),.ci(co1_14));
  fa u_csa2_15 (.s(sum2_15),.co(co2_15),.a(pp3_13),.b(sum1_16),.ci(co1_15));
  fa u_csa2_16 (.s(sum2_16),.co(co2_16),.a(pp3_14),.b(sum1_17),.ci(co1_16));
  fa u_csa2_17 (.s(sum2_17),.co(co2_17),.a(pp3_15),.b(sum1_18),.ci(co1_17));
  fa u_csa2_18 (.s(sum2_18),.co(co2_18),.a(pp3_16),.b(sum1_19),.ci(co1_18));
  fa u_csa2_19 (.s(sum2_19),.co(co2_19),.a(pp3_17),.b(sum1_20),.ci(co1_19));
  fa u_csa2_20 (.s(sum2_20),.co(co2_20),.a(pp3_18),.b(sum1_21),.ci(co1_20));
  fa u_csa2_21 (.s(sum2_21),.co(co2_21),.a(pp3_19),.b(sum1_22),.ci(co1_21));
  fa u_csa2_22 (.s(sum2_22),.co(co2_22),.a(pp3_20),.b(sum1_23),.ci(co1_22));
  fa u_csa2_23 (.s(sum2_23),.co(co2_23),.a(pp3_21),.b(sum1_24),.ci(co1_23));
  fa u_csa2_24 (.s(sum2_24),.co(co2_24),.a(pp3_22),.b(sum1_25),.ci(co1_24));
  fa u_csa2_25 (.s(sum2_25),.co(co2_25),.a(pp3_23),.b(sum1_26),.ci(co1_25));
  fa u_csa2_26 (.s(sum2_26),.co(co2_26),.a(pp3_24),.b(sum1_27),.ci(co1_26));
  fa u_csa2_27 (.s(sum2_27),.co(co2_27),.a(pp3_25),.b(sum1_28),.ci(co1_27));
  fa u_csa2_28 (.s(sum2_28),.co(co2_28),.a(pp3_26),.b(sum1_29),.ci(co1_28));
  fa u_csa2_29 (.s(sum2_29),.co(co2_29),.a(pp3_27),.b(sum1_30),.ci(co1_29));
  fa u_csa2_30 (.s(sum2_30),.co(co2_30),.a(pp3_28),.b(sum1_31),.ci(co1_30));
  fa u_csa2_31 (.s(sum2_31),.co(co2_31),.a(pp3_29),.b(sum1_32),.ci(co1_31));
  fa u_csa2_32 (.s(sum2_32),.co(co2_32),.a(pp3_30),.b(sum1_33),.ci(co1_32));
  fa u_csa2_33 (.s(sum2_33),.co(co2_33),.a(pp3_31),.b(sum1_34),.ci(co1_33));
  fa u_csa2_34 (.s(sum2_34),.co(co2_34),.a(pp3_32),.b(sum1_35),.ci(co1_34));
  fa u_csa2_35 (.s(sum2_35),.co(co2_35),.a(pp3_33),.b(sum1_36),.ci(co1_35));
  fa u_csa2_36 (.s(sum2_36),.co(co2_36),.a(pp3_34),.b(sum1_37),.ci(co1_36));
  assign sum2_37=pp3_35;
  assign co2_37=sig0;
  assign sum2_38=pp3_36;
  //CSA Row 3 
  ha u_csa3_0 (.s(sum3_0),.co(co3_0),.a(sum2_1),.b(co2_0));
  ha u_csa3_1 (.s(sum3_1),.co(co3_1),.a(sum2_2),.b(co2_1));
  ha u_csa3_2 (.s(sum3_2),.co(co3_2),.a(sum2_3),.b(co2_2));
  fa u_csa3_3 (.s(sum3_3),.co(co3_3),.a(pp4_0),.b(sum2_4),.ci(co2_3));
  fa u_csa3_4 (.s(sum3_4),.co(co3_4),.a(pp4_1),.b(sum2_5),.ci(co2_4));
  fa u_csa3_5 (.s(sum3_5),.co(co3_5),.a(pp4_2),.b(sum2_6),.ci(co2_5));
  fa u_csa3_6 (.s(sum3_6),.co(co3_6),.a(pp4_3),.b(sum2_7),.ci(co2_6));
  fa u_csa3_7 (.s(sum3_7),.co(co3_7),.a(pp4_4),.b(sum2_8),.ci(co2_7));
  fa u_csa3_8 (.s(sum3_8),.co(co3_8),.a(pp4_5),.b(sum2_9),.ci(co2_8));
  fa u_csa3_9 (.s(sum3_9),.co(co3_9),.a(pp4_6),.b(sum2_10),.ci(co2_9));
  fa u_csa3_10 (.s(sum3_10),.co(co3_10),.a(pp4_7),.b(sum2_11),.ci(co2_10));
  fa u_csa3_11 (.s(sum3_11),.co(co3_11),.a(pp4_8),.b(sum2_12),.ci(co2_11));
  fa u_csa3_12 (.s(sum3_12),.co(co3_12),.a(pp4_9),.b(sum2_13),.ci(co2_12));
  fa u_csa3_13 (.s(sum3_13),.co(co3_13),.a(pp4_10),.b(sum2_14),.ci(co2_13));
  fa u_csa3_14 (.s(sum3_14),.co(co3_14),.a(pp4_11),.b(sum2_15),.ci(co2_14));
  fa u_csa3_15 (.s(sum3_15),.co(co3_15),.a(pp4_12),.b(sum2_16),.ci(co2_15));
  fa u_csa3_16 (.s(sum3_16),.co(co3_16),.a(pp4_13),.b(sum2_17),.ci(co2_16));
  fa u_csa3_17 (.s(sum3_17),.co(co3_17),.a(pp4_14),.b(sum2_18),.ci(co2_17));
  fa u_csa3_18 (.s(sum3_18),.co(co3_18),.a(pp4_15),.b(sum2_19),.ci(co2_18));
  fa u_csa3_19 (.s(sum3_19),.co(co3_19),.a(pp4_16),.b(sum2_20),.ci(co2_19));
  fa u_csa3_20 (.s(sum3_20),.co(co3_20),.a(pp4_17),.b(sum2_21),.ci(co2_20));
  fa u_csa3_21 (.s(sum3_21),.co(co3_21),.a(pp4_18),.b(sum2_22),.ci(co2_21));
  fa u_csa3_22 (.s(sum3_22),.co(co3_22),.a(pp4_19),.b(sum2_23),.ci(co2_22));
  fa u_csa3_23 (.s(sum3_23),.co(co3_23),.a(pp4_20),.b(sum2_24),.ci(co2_23));
  fa u_csa3_24 (.s(sum3_24),.co(co3_24),.a(pp4_21),.b(sum2_25),.ci(co2_24));
  fa u_csa3_25 (.s(sum3_25),.co(co3_25),.a(pp4_22),.b(sum2_26),.ci(co2_25));
  fa u_csa3_26 (.s(sum3_26),.co(co3_26),.a(pp4_23),.b(sum2_27),.ci(co2_26));
  fa u_csa3_27 (.s(sum3_27),.co(co3_27),.a(pp4_24),.b(sum2_28),.ci(co2_27));
  fa u_csa3_28 (.s(sum3_28),.co(co3_28),.a(pp4_25),.b(sum2_29),.ci(co2_28));
  fa u_csa3_29 (.s(sum3_29),.co(co3_29),.a(pp4_26),.b(sum2_30),.ci(co2_29));
  fa u_csa3_30 (.s(sum3_30),.co(co3_30),.a(pp4_27),.b(sum2_31),.ci(co2_30));
  fa u_csa3_31 (.s(sum3_31),.co(co3_31),.a(pp4_28),.b(sum2_32),.ci(co2_31));
  fa u_csa3_32 (.s(sum3_32),.co(co3_32),.a(pp4_29),.b(sum2_33),.ci(co2_32));
  fa u_csa3_33 (.s(sum3_33),.co(co3_33),.a(pp4_30),.b(sum2_34),.ci(co2_33));
  fa u_csa3_34 (.s(sum3_34),.co(co3_34),.a(pp4_31),.b(sum2_35),.ci(co2_34));
  fa u_csa3_35 (.s(sum3_35),.co(co3_35),.a(pp4_32),.b(sum2_36),.ci(co2_35));
  fa u_csa3_36 (.s(sum3_36),.co(co3_36),.a(pp4_33),.b(sum2_37),.ci(co2_36));
  fa u_csa3_37 (.s(sum3_37),.co(co3_37),.a(pp4_34),.b(sum2_38),.ci(co2_37));
  assign sum3_38=pp4_35;
  assign co3_38=sig0;
  assign sum3_39=pp4_36;
  //CSA Row 4 
  ha u_csa4_0 (.s(sum4_0),.co(co4_0),.a(sum3_1),.b(co3_0));
  ha u_csa4_1 (.s(sum4_1),.co(co4_1),.a(sum3_2),.b(co3_1));
  ha u_csa4_2 (.s(sum4_2),.co(co4_2),.a(sum3_3),.b(co3_2));
  ha u_csa4_3 (.s(sum4_3),.co(co4_3),.a(sum3_4),.b(co3_3));
  fa u_csa4_4 (.s(sum4_4),.co(co4_4),.a(pp5_0),.b(sum3_5),.ci(co3_4));
  fa u_csa4_5 (.s(sum4_5),.co(co4_5),.a(pp5_1),.b(sum3_6),.ci(co3_5));
  fa u_csa4_6 (.s(sum4_6),.co(co4_6),.a(pp5_2),.b(sum3_7),.ci(co3_6));
  fa u_csa4_7 (.s(sum4_7),.co(co4_7),.a(pp5_3),.b(sum3_8),.ci(co3_7));
  fa u_csa4_8 (.s(sum4_8),.co(co4_8),.a(pp5_4),.b(sum3_9),.ci(co3_8));
  fa u_csa4_9 (.s(sum4_9),.co(co4_9),.a(pp5_5),.b(sum3_10),.ci(co3_9));
  fa u_csa4_10 (.s(sum4_10),.co(co4_10),.a(pp5_6),.b(sum3_11),.ci(co3_10));
  fa u_csa4_11 (.s(sum4_11),.co(co4_11),.a(pp5_7),.b(sum3_12),.ci(co3_11));
  fa u_csa4_12 (.s(sum4_12),.co(co4_12),.a(pp5_8),.b(sum3_13),.ci(co3_12));
  fa u_csa4_13 (.s(sum4_13),.co(co4_13),.a(pp5_9),.b(sum3_14),.ci(co3_13));
  fa u_csa4_14 (.s(sum4_14),.co(co4_14),.a(pp5_10),.b(sum3_15),.ci(co3_14));
  fa u_csa4_15 (.s(sum4_15),.co(co4_15),.a(pp5_11),.b(sum3_16),.ci(co3_15));
  fa u_csa4_16 (.s(sum4_16),.co(co4_16),.a(pp5_12),.b(sum3_17),.ci(co3_16));
  fa u_csa4_17 (.s(sum4_17),.co(co4_17),.a(pp5_13),.b(sum3_18),.ci(co3_17));
  fa u_csa4_18 (.s(sum4_18),.co(co4_18),.a(pp5_14),.b(sum3_19),.ci(co3_18));
  fa u_csa4_19 (.s(sum4_19),.co(co4_19),.a(pp5_15),.b(sum3_20),.ci(co3_19));
  fa u_csa4_20 (.s(sum4_20),.co(co4_20),.a(pp5_16),.b(sum3_21),.ci(co3_20));
  fa u_csa4_21 (.s(sum4_21),.co(co4_21),.a(pp5_17),.b(sum3_22),.ci(co3_21));
  fa u_csa4_22 (.s(sum4_22),.co(co4_22),.a(pp5_18),.b(sum3_23),.ci(co3_22));
  fa u_csa4_23 (.s(sum4_23),.co(co4_23),.a(pp5_19),.b(sum3_24),.ci(co3_23));
  fa u_csa4_24 (.s(sum4_24),.co(co4_24),.a(pp5_20),.b(sum3_25),.ci(co3_24));
  fa u_csa4_25 (.s(sum4_25),.co(co4_25),.a(pp5_21),.b(sum3_26),.ci(co3_25));
  fa u_csa4_26 (.s(sum4_26),.co(co4_26),.a(pp5_22),.b(sum3_27),.ci(co3_26));
  fa u_csa4_27 (.s(sum4_27),.co(co4_27),.a(pp5_23),.b(sum3_28),.ci(co3_27));
  fa u_csa4_28 (.s(sum4_28),.co(co4_28),.a(pp5_24),.b(sum3_29),.ci(co3_28));
  fa u_csa4_29 (.s(sum4_29),.co(co4_29),.a(pp5_25),.b(sum3_30),.ci(co3_29));
  fa u_csa4_30 (.s(sum4_30),.co(co4_30),.a(pp5_26),.b(sum3_31),.ci(co3_30));
  fa u_csa4_31 (.s(sum4_31),.co(co4_31),.a(pp5_27),.b(sum3_32),.ci(co3_31));
  fa u_csa4_32 (.s(sum4_32),.co(co4_32),.a(pp5_28),.b(sum3_33),.ci(co3_32));
  fa u_csa4_33 (.s(sum4_33),.co(co4_33),.a(pp5_29),.b(sum3_34),.ci(co3_33));
  fa u_csa4_34 (.s(sum4_34),.co(co4_34),.a(pp5_30),.b(sum3_35),.ci(co3_34));
  fa u_csa4_35 (.s(sum4_35),.co(co4_35),.a(pp5_31),.b(sum3_36),.ci(co3_35));
  fa u_csa4_36 (.s(sum4_36),.co(co4_36),.a(pp5_32),.b(sum3_37),.ci(co3_36));
  fa u_csa4_37 (.s(sum4_37),.co(co4_37),.a(pp5_33),.b(sum3_38),.ci(co3_37));
  fa u_csa4_38 (.s(sum4_38),.co(co4_38),.a(pp5_34),.b(sum3_39),.ci(co3_38));
  assign sum4_39=pp5_35;
  assign co4_39=sig0;
  assign sum4_40=pp5_36;
  //CSA Row 5 
  ha u_csa5_0 (.s(sum5_0),.co(co5_0),.a(sum4_1),.b(co4_0));
  ha u_csa5_1 (.s(sum5_1),.co(co5_1),.a(sum4_2),.b(co4_1));
  ha u_csa5_2 (.s(sum5_2),.co(co5_2),.a(sum4_3),.b(co4_2));
  ha u_csa5_3 (.s(sum5_3),.co(co5_3),.a(sum4_4),.b(co4_3));
  ha u_csa5_4 (.s(sum5_4),.co(co5_4),.a(sum4_5),.b(co4_4));
  fa u_csa5_5 (.s(sum5_5),.co(co5_5),.a(pp6_0),.b(sum4_6),.ci(co4_5));
  fa u_csa5_6 (.s(sum5_6),.co(co5_6),.a(pp6_1),.b(sum4_7),.ci(co4_6));
  fa u_csa5_7 (.s(sum5_7),.co(co5_7),.a(pp6_2),.b(sum4_8),.ci(co4_7));
  fa u_csa5_8 (.s(sum5_8),.co(co5_8),.a(pp6_3),.b(sum4_9),.ci(co4_8));
  fa u_csa5_9 (.s(sum5_9),.co(co5_9),.a(pp6_4),.b(sum4_10),.ci(co4_9));
  fa u_csa5_10 (.s(sum5_10),.co(co5_10),.a(pp6_5),.b(sum4_11),.ci(co4_10));
  fa u_csa5_11 (.s(sum5_11),.co(co5_11),.a(pp6_6),.b(sum4_12),.ci(co4_11));
  fa u_csa5_12 (.s(sum5_12),.co(co5_12),.a(pp6_7),.b(sum4_13),.ci(co4_12));
  fa u_csa5_13 (.s(sum5_13),.co(co5_13),.a(pp6_8),.b(sum4_14),.ci(co4_13));
  fa u_csa5_14 (.s(sum5_14),.co(co5_14),.a(pp6_9),.b(sum4_15),.ci(co4_14));
  fa u_csa5_15 (.s(sum5_15),.co(co5_15),.a(pp6_10),.b(sum4_16),.ci(co4_15));
  fa u_csa5_16 (.s(sum5_16),.co(co5_16),.a(pp6_11),.b(sum4_17),.ci(co4_16));
  fa u_csa5_17 (.s(sum5_17),.co(co5_17),.a(pp6_12),.b(sum4_18),.ci(co4_17));
  fa u_csa5_18 (.s(sum5_18),.co(co5_18),.a(pp6_13),.b(sum4_19),.ci(co4_18));
  fa u_csa5_19 (.s(sum5_19),.co(co5_19),.a(pp6_14),.b(sum4_20),.ci(co4_19));
  fa u_csa5_20 (.s(sum5_20),.co(co5_20),.a(pp6_15),.b(sum4_21),.ci(co4_20));
  fa u_csa5_21 (.s(sum5_21),.co(co5_21),.a(pp6_16),.b(sum4_22),.ci(co4_21));
  fa u_csa5_22 (.s(sum5_22),.co(co5_22),.a(pp6_17),.b(sum4_23),.ci(co4_22));
  fa u_csa5_23 (.s(sum5_23),.co(co5_23),.a(pp6_18),.b(sum4_24),.ci(co4_23));
  fa u_csa5_24 (.s(sum5_24),.co(co5_24),.a(pp6_19),.b(sum4_25),.ci(co4_24));
  fa u_csa5_25 (.s(sum5_25),.co(co5_25),.a(pp6_20),.b(sum4_26),.ci(co4_25));
  fa u_csa5_26 (.s(sum5_26),.co(co5_26),.a(pp6_21),.b(sum4_27),.ci(co4_26));
  fa u_csa5_27 (.s(sum5_27),.co(co5_27),.a(pp6_22),.b(sum4_28),.ci(co4_27));
  fa u_csa5_28 (.s(sum5_28),.co(co5_28),.a(pp6_23),.b(sum4_29),.ci(co4_28));
  fa u_csa5_29 (.s(sum5_29),.co(co5_29),.a(pp6_24),.b(sum4_30),.ci(co4_29));
  fa u_csa5_30 (.s(sum5_30),.co(co5_30),.a(pp6_25),.b(sum4_31),.ci(co4_30));
  fa u_csa5_31 (.s(sum5_31),.co(co5_31),.a(pp6_26),.b(sum4_32),.ci(co4_31));
  fa u_csa5_32 (.s(sum5_32),.co(co5_32),.a(pp6_27),.b(sum4_33),.ci(co4_32));
  fa u_csa5_33 (.s(sum5_33),.co(co5_33),.a(pp6_28),.b(sum4_34),.ci(co4_33));
  fa u_csa5_34 (.s(sum5_34),.co(co5_34),.a(pp6_29),.b(sum4_35),.ci(co4_34));
  fa u_csa5_35 (.s(sum5_35),.co(co5_35),.a(pp6_30),.b(sum4_36),.ci(co4_35));
  fa u_csa5_36 (.s(sum5_36),.co(co5_36),.a(pp6_31),.b(sum4_37),.ci(co4_36));
  fa u_csa5_37 (.s(sum5_37),.co(co5_37),.a(pp6_32),.b(sum4_38),.ci(co4_37));
  fa u_csa5_38 (.s(sum5_38),.co(co5_38),.a(pp6_33),.b(sum4_39),.ci(co4_38));
  fa u_csa5_39 (.s(sum5_39),.co(co5_39),.a(pp6_34),.b(sum4_40),.ci(co4_39));
  assign sum5_40=pp6_35;
  assign co5_40=sig0;
  assign sum5_41=pp6_36;
  //CSA Row 6 
  ha u_csa6_0 (.s(sum6_0),.co(co6_0),.a(sum5_1),.b(co5_0));
  ha u_csa6_1 (.s(sum6_1),.co(co6_1),.a(sum5_2),.b(co5_1));
  ha u_csa6_2 (.s(sum6_2),.co(co6_2),.a(sum5_3),.b(co5_2));
  ha u_csa6_3 (.s(sum6_3),.co(co6_3),.a(sum5_4),.b(co5_3));
  ha u_csa6_4 (.s(sum6_4),.co(co6_4),.a(sum5_5),.b(co5_4));
  ha u_csa6_5 (.s(sum6_5),.co(co6_5),.a(sum5_6),.b(co5_5));
  fa u_csa6_6 (.s(sum6_6),.co(co6_6),.a(pp7_0),.b(sum5_7),.ci(co5_6));
  fa u_csa6_7 (.s(sum6_7),.co(co6_7),.a(pp7_1),.b(sum5_8),.ci(co5_7));
  fa u_csa6_8 (.s(sum6_8),.co(co6_8),.a(pp7_2),.b(sum5_9),.ci(co5_8));
  fa u_csa6_9 (.s(sum6_9),.co(co6_9),.a(pp7_3),.b(sum5_10),.ci(co5_9));
  fa u_csa6_10 (.s(sum6_10),.co(co6_10),.a(pp7_4),.b(sum5_11),.ci(co5_10));
  fa u_csa6_11 (.s(sum6_11),.co(co6_11),.a(pp7_5),.b(sum5_12),.ci(co5_11));
  fa u_csa6_12 (.s(sum6_12),.co(co6_12),.a(pp7_6),.b(sum5_13),.ci(co5_12));
  fa u_csa6_13 (.s(sum6_13),.co(co6_13),.a(pp7_7),.b(sum5_14),.ci(co5_13));
  fa u_csa6_14 (.s(sum6_14),.co(co6_14),.a(pp7_8),.b(sum5_15),.ci(co5_14));
  fa u_csa6_15 (.s(sum6_15),.co(co6_15),.a(pp7_9),.b(sum5_16),.ci(co5_15));
  fa u_csa6_16 (.s(sum6_16),.co(co6_16),.a(pp7_10),.b(sum5_17),.ci(co5_16));
  fa u_csa6_17 (.s(sum6_17),.co(co6_17),.a(pp7_11),.b(sum5_18),.ci(co5_17));
  fa u_csa6_18 (.s(sum6_18),.co(co6_18),.a(pp7_12),.b(sum5_19),.ci(co5_18));
  fa u_csa6_19 (.s(sum6_19),.co(co6_19),.a(pp7_13),.b(sum5_20),.ci(co5_19));
  fa u_csa6_20 (.s(sum6_20),.co(co6_20),.a(pp7_14),.b(sum5_21),.ci(co5_20));
  fa u_csa6_21 (.s(sum6_21),.co(co6_21),.a(pp7_15),.b(sum5_22),.ci(co5_21));
  fa u_csa6_22 (.s(sum6_22),.co(co6_22),.a(pp7_16),.b(sum5_23),.ci(co5_22));
  fa u_csa6_23 (.s(sum6_23),.co(co6_23),.a(pp7_17),.b(sum5_24),.ci(co5_23));
  fa u_csa6_24 (.s(sum6_24),.co(co6_24),.a(pp7_18),.b(sum5_25),.ci(co5_24));
  fa u_csa6_25 (.s(sum6_25),.co(co6_25),.a(pp7_19),.b(sum5_26),.ci(co5_25));
  fa u_csa6_26 (.s(sum6_26),.co(co6_26),.a(pp7_20),.b(sum5_27),.ci(co5_26));
  fa u_csa6_27 (.s(sum6_27),.co(co6_27),.a(pp7_21),.b(sum5_28),.ci(co5_27));
  fa u_csa6_28 (.s(sum6_28),.co(co6_28),.a(pp7_22),.b(sum5_29),.ci(co5_28));
  fa u_csa6_29 (.s(sum6_29),.co(co6_29),.a(pp7_23),.b(sum5_30),.ci(co5_29));
  fa u_csa6_30 (.s(sum6_30),.co(co6_30),.a(pp7_24),.b(sum5_31),.ci(co5_30));
  fa u_csa6_31 (.s(sum6_31),.co(co6_31),.a(pp7_25),.b(sum5_32),.ci(co5_31));
  fa u_csa6_32 (.s(sum6_32),.co(co6_32),.a(pp7_26),.b(sum5_33),.ci(co5_32));
  fa u_csa6_33 (.s(sum6_33),.co(co6_33),.a(pp7_27),.b(sum5_34),.ci(co5_33));
  fa u_csa6_34 (.s(sum6_34),.co(co6_34),.a(pp7_28),.b(sum5_35),.ci(co5_34));
  fa u_csa6_35 (.s(sum6_35),.co(co6_35),.a(pp7_29),.b(sum5_36),.ci(co5_35));
  fa u_csa6_36 (.s(sum6_36),.co(co6_36),.a(pp7_30),.b(sum5_37),.ci(co5_36));
  fa u_csa6_37 (.s(sum6_37),.co(co6_37),.a(pp7_31),.b(sum5_38),.ci(co5_37));
  fa u_csa6_38 (.s(sum6_38),.co(co6_38),.a(pp7_32),.b(sum5_39),.ci(co5_38));
  fa u_csa6_39 (.s(sum6_39),.co(co6_39),.a(pp7_33),.b(sum5_40),.ci(co5_39));
  fa u_csa6_40 (.s(sum6_40),.co(co6_40),.a(pp7_34),.b(sum5_41),.ci(co5_40));
  assign sum6_41=pp7_35;
  assign co6_41=sig0;
  assign sum6_42=pp7_36;
  //CSA Row 7 
  ha u_csa7_0 (.s(sum7_0),.co(co7_0),.a(sum6_1),.b(co6_0));
  ha u_csa7_1 (.s(sum7_1),.co(co7_1),.a(sum6_2),.b(co6_1));
  ha u_csa7_2 (.s(sum7_2),.co(co7_2),.a(sum6_3),.b(co6_2));
  ha u_csa7_3 (.s(sum7_3),.co(co7_3),.a(sum6_4),.b(co6_3));
  ha u_csa7_4 (.s(sum7_4),.co(co7_4),.a(sum6_5),.b(co6_4));
  ha u_csa7_5 (.s(sum7_5),.co(co7_5),.a(sum6_6),.b(co6_5));
  ha u_csa7_6 (.s(sum7_6),.co(co7_6),.a(sum6_7),.b(co6_6));
  fa u_csa7_7 (.s(sum7_7),.co(co7_7),.a(pp8_0),.b(sum6_8),.ci(co6_7));
  fa u_csa7_8 (.s(sum7_8),.co(co7_8),.a(pp8_1),.b(sum6_9),.ci(co6_8));
  fa u_csa7_9 (.s(sum7_9),.co(co7_9),.a(pp8_2),.b(sum6_10),.ci(co6_9));
  fa u_csa7_10 (.s(sum7_10),.co(co7_10),.a(pp8_3),.b(sum6_11),.ci(co6_10));
  fa u_csa7_11 (.s(sum7_11),.co(co7_11),.a(pp8_4),.b(sum6_12),.ci(co6_11));
  fa u_csa7_12 (.s(sum7_12),.co(co7_12),.a(pp8_5),.b(sum6_13),.ci(co6_12));
  fa u_csa7_13 (.s(sum7_13),.co(co7_13),.a(pp8_6),.b(sum6_14),.ci(co6_13));
  fa u_csa7_14 (.s(sum7_14),.co(co7_14),.a(pp8_7),.b(sum6_15),.ci(co6_14));
  fa u_csa7_15 (.s(sum7_15),.co(co7_15),.a(pp8_8),.b(sum6_16),.ci(co6_15));
  fa u_csa7_16 (.s(sum7_16),.co(co7_16),.a(pp8_9),.b(sum6_17),.ci(co6_16));
  fa u_csa7_17 (.s(sum7_17),.co(co7_17),.a(pp8_10),.b(sum6_18),.ci(co6_17));
  fa u_csa7_18 (.s(sum7_18),.co(co7_18),.a(pp8_11),.b(sum6_19),.ci(co6_18));
  fa u_csa7_19 (.s(sum7_19),.co(co7_19),.a(pp8_12),.b(sum6_20),.ci(co6_19));
  fa u_csa7_20 (.s(sum7_20),.co(co7_20),.a(pp8_13),.b(sum6_21),.ci(co6_20));
  fa u_csa7_21 (.s(sum7_21),.co(co7_21),.a(pp8_14),.b(sum6_22),.ci(co6_21));
  fa u_csa7_22 (.s(sum7_22),.co(co7_22),.a(pp8_15),.b(sum6_23),.ci(co6_22));
  fa u_csa7_23 (.s(sum7_23),.co(co7_23),.a(pp8_16),.b(sum6_24),.ci(co6_23));
  fa u_csa7_24 (.s(sum7_24),.co(co7_24),.a(pp8_17),.b(sum6_25),.ci(co6_24));
  fa u_csa7_25 (.s(sum7_25),.co(co7_25),.a(pp8_18),.b(sum6_26),.ci(co6_25));
  fa u_csa7_26 (.s(sum7_26),.co(co7_26),.a(pp8_19),.b(sum6_27),.ci(co6_26));
  fa u_csa7_27 (.s(sum7_27),.co(co7_27),.a(pp8_20),.b(sum6_28),.ci(co6_27));
  fa u_csa7_28 (.s(sum7_28),.co(co7_28),.a(pp8_21),.b(sum6_29),.ci(co6_28));
  fa u_csa7_29 (.s(sum7_29),.co(co7_29),.a(pp8_22),.b(sum6_30),.ci(co6_29));
  fa u_csa7_30 (.s(sum7_30),.co(co7_30),.a(pp8_23),.b(sum6_31),.ci(co6_30));
  fa u_csa7_31 (.s(sum7_31),.co(co7_31),.a(pp8_24),.b(sum6_32),.ci(co6_31));
  fa u_csa7_32 (.s(sum7_32),.co(co7_32),.a(pp8_25),.b(sum6_33),.ci(co6_32));
  fa u_csa7_33 (.s(sum7_33),.co(co7_33),.a(pp8_26),.b(sum6_34),.ci(co6_33));
  fa u_csa7_34 (.s(sum7_34),.co(co7_34),.a(pp8_27),.b(sum6_35),.ci(co6_34));
  fa u_csa7_35 (.s(sum7_35),.co(co7_35),.a(pp8_28),.b(sum6_36),.ci(co6_35));
  fa u_csa7_36 (.s(sum7_36),.co(co7_36),.a(pp8_29),.b(sum6_37),.ci(co6_36));
  fa u_csa7_37 (.s(sum7_37),.co(co7_37),.a(pp8_30),.b(sum6_38),.ci(co6_37));
  fa u_csa7_38 (.s(sum7_38),.co(co7_38),.a(pp8_31),.b(sum6_39),.ci(co6_38));
  fa u_csa7_39 (.s(sum7_39),.co(co7_39),.a(pp8_32),.b(sum6_40),.ci(co6_39));
  fa u_csa7_40 (.s(sum7_40),.co(co7_40),.a(pp8_33),.b(sum6_41),.ci(co6_40));
  fa u_csa7_41 (.s(sum7_41),.co(co7_41),.a(pp8_34),.b(sum6_42),.ci(co6_41));
  assign sum7_42=pp8_35;
  assign co7_42=sig0;
  assign sum7_43=pp8_36;
  //CSA Row 8 
  ha u_csa8_0 (.s(sum8_0),.co(co8_0),.a(sum7_1),.b(co7_0));
  ha u_csa8_1 (.s(sum8_1),.co(co8_1),.a(sum7_2),.b(co7_1));
  ha u_csa8_2 (.s(sum8_2),.co(co8_2),.a(sum7_3),.b(co7_2));
  ha u_csa8_3 (.s(sum8_3),.co(co8_3),.a(sum7_4),.b(co7_3));
  ha u_csa8_4 (.s(sum8_4),.co(co8_4),.a(sum7_5),.b(co7_4));
  ha u_csa8_5 (.s(sum8_5),.co(co8_5),.a(sum7_6),.b(co7_5));
  ha u_csa8_6 (.s(sum8_6),.co(co8_6),.a(sum7_7),.b(co7_6));
  ha u_csa8_7 (.s(sum8_7),.co(co8_7),.a(sum7_8),.b(co7_7));
  fa u_csa8_8 (.s(sum8_8),.co(co8_8),.a(pp9_0),.b(sum7_9),.ci(co7_8));
  fa u_csa8_9 (.s(sum8_9),.co(co8_9),.a(pp9_1),.b(sum7_10),.ci(co7_9));
  fa u_csa8_10 (.s(sum8_10),.co(co8_10),.a(pp9_2),.b(sum7_11),.ci(co7_10));
  fa u_csa8_11 (.s(sum8_11),.co(co8_11),.a(pp9_3),.b(sum7_12),.ci(co7_11));
  fa u_csa8_12 (.s(sum8_12),.co(co8_12),.a(pp9_4),.b(sum7_13),.ci(co7_12));
  fa u_csa8_13 (.s(sum8_13),.co(co8_13),.a(pp9_5),.b(sum7_14),.ci(co7_13));
  fa u_csa8_14 (.s(sum8_14),.co(co8_14),.a(pp9_6),.b(sum7_15),.ci(co7_14));
  fa u_csa8_15 (.s(sum8_15),.co(co8_15),.a(pp9_7),.b(sum7_16),.ci(co7_15));
  fa u_csa8_16 (.s(sum8_16),.co(co8_16),.a(pp9_8),.b(sum7_17),.ci(co7_16));
  fa u_csa8_17 (.s(sum8_17),.co(co8_17),.a(pp9_9),.b(sum7_18),.ci(co7_17));
  fa u_csa8_18 (.s(sum8_18),.co(co8_18),.a(pp9_10),.b(sum7_19),.ci(co7_18));
  fa u_csa8_19 (.s(sum8_19),.co(co8_19),.a(pp9_11),.b(sum7_20),.ci(co7_19));
  fa u_csa8_20 (.s(sum8_20),.co(co8_20),.a(pp9_12),.b(sum7_21),.ci(co7_20));
  fa u_csa8_21 (.s(sum8_21),.co(co8_21),.a(pp9_13),.b(sum7_22),.ci(co7_21));
  fa u_csa8_22 (.s(sum8_22),.co(co8_22),.a(pp9_14),.b(sum7_23),.ci(co7_22));
  fa u_csa8_23 (.s(sum8_23),.co(co8_23),.a(pp9_15),.b(sum7_24),.ci(co7_23));
  fa u_csa8_24 (.s(sum8_24),.co(co8_24),.a(pp9_16),.b(sum7_25),.ci(co7_24));
  fa u_csa8_25 (.s(sum8_25),.co(co8_25),.a(pp9_17),.b(sum7_26),.ci(co7_25));
  fa u_csa8_26 (.s(sum8_26),.co(co8_26),.a(pp9_18),.b(sum7_27),.ci(co7_26));
  fa u_csa8_27 (.s(sum8_27),.co(co8_27),.a(pp9_19),.b(sum7_28),.ci(co7_27));
  fa u_csa8_28 (.s(sum8_28),.co(co8_28),.a(pp9_20),.b(sum7_29),.ci(co7_28));
  fa u_csa8_29 (.s(sum8_29),.co(co8_29),.a(pp9_21),.b(sum7_30),.ci(co7_29));
  fa u_csa8_30 (.s(sum8_30),.co(co8_30),.a(pp9_22),.b(sum7_31),.ci(co7_30));
  fa u_csa8_31 (.s(sum8_31),.co(co8_31),.a(pp9_23),.b(sum7_32),.ci(co7_31));
  fa u_csa8_32 (.s(sum8_32),.co(co8_32),.a(pp9_24),.b(sum7_33),.ci(co7_32));
  fa u_csa8_33 (.s(sum8_33),.co(co8_33),.a(pp9_25),.b(sum7_34),.ci(co7_33));
  fa u_csa8_34 (.s(sum8_34),.co(co8_34),.a(pp9_26),.b(sum7_35),.ci(co7_34));
  fa u_csa8_35 (.s(sum8_35),.co(co8_35),.a(pp9_27),.b(sum7_36),.ci(co7_35));
  fa u_csa8_36 (.s(sum8_36),.co(co8_36),.a(pp9_28),.b(sum7_37),.ci(co7_36));
  fa u_csa8_37 (.s(sum8_37),.co(co8_37),.a(pp9_29),.b(sum7_38),.ci(co7_37));
  fa u_csa8_38 (.s(sum8_38),.co(co8_38),.a(pp9_30),.b(sum7_39),.ci(co7_38));
  fa u_csa8_39 (.s(sum8_39),.co(co8_39),.a(pp9_31),.b(sum7_40),.ci(co7_39));
  fa u_csa8_40 (.s(sum8_40),.co(co8_40),.a(pp9_32),.b(sum7_41),.ci(co7_40));
  fa u_csa8_41 (.s(sum8_41),.co(co8_41),.a(pp9_33),.b(sum7_42),.ci(co7_41));
  fa u_csa8_42 (.s(sum8_42),.co(co8_42),.a(pp9_34),.b(sum7_43),.ci(co7_42));
  assign sum8_43=pp9_35;
  assign co8_43=sig0;
  assign sum8_44=pp9_36;
  //CSA Row 9 
  ha u_csa9_0 (.s(sum9_0),.co(co9_0),.a(sum8_1),.b(co8_0));
  ha u_csa9_1 (.s(sum9_1),.co(co9_1),.a(sum8_2),.b(co8_1));
  ha u_csa9_2 (.s(sum9_2),.co(co9_2),.a(sum8_3),.b(co8_2));
  ha u_csa9_3 (.s(sum9_3),.co(co9_3),.a(sum8_4),.b(co8_3));
  ha u_csa9_4 (.s(sum9_4),.co(co9_4),.a(sum8_5),.b(co8_4));
  ha u_csa9_5 (.s(sum9_5),.co(co9_5),.a(sum8_6),.b(co8_5));
  ha u_csa9_6 (.s(sum9_6),.co(co9_6),.a(sum8_7),.b(co8_6));
  ha u_csa9_7 (.s(sum9_7),.co(co9_7),.a(sum8_8),.b(co8_7));
  ha u_csa9_8 (.s(sum9_8),.co(co9_8),.a(sum8_9),.b(co8_8));
  fa u_csa9_9 (.s(sum9_9),.co(co9_9),.a(pp10_0),.b(sum8_10),.ci(co8_9));
  fa u_csa9_10 (.s(sum9_10),.co(co9_10),.a(pp10_1),.b(sum8_11),.ci(co8_10));
  fa u_csa9_11 (.s(sum9_11),.co(co9_11),.a(pp10_2),.b(sum8_12),.ci(co8_11));
  fa u_csa9_12 (.s(sum9_12),.co(co9_12),.a(pp10_3),.b(sum8_13),.ci(co8_12));
  fa u_csa9_13 (.s(sum9_13),.co(co9_13),.a(pp10_4),.b(sum8_14),.ci(co8_13));
  fa u_csa9_14 (.s(sum9_14),.co(co9_14),.a(pp10_5),.b(sum8_15),.ci(co8_14));
  fa u_csa9_15 (.s(sum9_15),.co(co9_15),.a(pp10_6),.b(sum8_16),.ci(co8_15));
  fa u_csa9_16 (.s(sum9_16),.co(co9_16),.a(pp10_7),.b(sum8_17),.ci(co8_16));
  fa u_csa9_17 (.s(sum9_17),.co(co9_17),.a(pp10_8),.b(sum8_18),.ci(co8_17));
  fa u_csa9_18 (.s(sum9_18),.co(co9_18),.a(pp10_9),.b(sum8_19),.ci(co8_18));
  fa u_csa9_19 (.s(sum9_19),.co(co9_19),.a(pp10_10),.b(sum8_20),.ci(co8_19));
  fa u_csa9_20 (.s(sum9_20),.co(co9_20),.a(pp10_11),.b(sum8_21),.ci(co8_20));
  fa u_csa9_21 (.s(sum9_21),.co(co9_21),.a(pp10_12),.b(sum8_22),.ci(co8_21));
  fa u_csa9_22 (.s(sum9_22),.co(co9_22),.a(pp10_13),.b(sum8_23),.ci(co8_22));
  fa u_csa9_23 (.s(sum9_23),.co(co9_23),.a(pp10_14),.b(sum8_24),.ci(co8_23));
  fa u_csa9_24 (.s(sum9_24),.co(co9_24),.a(pp10_15),.b(sum8_25),.ci(co8_24));
  fa u_csa9_25 (.s(sum9_25),.co(co9_25),.a(pp10_16),.b(sum8_26),.ci(co8_25));
  fa u_csa9_26 (.s(sum9_26),.co(co9_26),.a(pp10_17),.b(sum8_27),.ci(co8_26));
  fa u_csa9_27 (.s(sum9_27),.co(co9_27),.a(pp10_18),.b(sum8_28),.ci(co8_27));
  fa u_csa9_28 (.s(sum9_28),.co(co9_28),.a(pp10_19),.b(sum8_29),.ci(co8_28));
  fa u_csa9_29 (.s(sum9_29),.co(co9_29),.a(pp10_20),.b(sum8_30),.ci(co8_29));
  fa u_csa9_30 (.s(sum9_30),.co(co9_30),.a(pp10_21),.b(sum8_31),.ci(co8_30));
  fa u_csa9_31 (.s(sum9_31),.co(co9_31),.a(pp10_22),.b(sum8_32),.ci(co8_31));
  fa u_csa9_32 (.s(sum9_32),.co(co9_32),.a(pp10_23),.b(sum8_33),.ci(co8_32));
  fa u_csa9_33 (.s(sum9_33),.co(co9_33),.a(pp10_24),.b(sum8_34),.ci(co8_33));
  fa u_csa9_34 (.s(sum9_34),.co(co9_34),.a(pp10_25),.b(sum8_35),.ci(co8_34));
  fa u_csa9_35 (.s(sum9_35),.co(co9_35),.a(pp10_26),.b(sum8_36),.ci(co8_35));
  fa u_csa9_36 (.s(sum9_36),.co(co9_36),.a(pp10_27),.b(sum8_37),.ci(co8_36));
  fa u_csa9_37 (.s(sum9_37),.co(co9_37),.a(pp10_28),.b(sum8_38),.ci(co8_37));
  fa u_csa9_38 (.s(sum9_38),.co(co9_38),.a(pp10_29),.b(sum8_39),.ci(co8_38));
  fa u_csa9_39 (.s(sum9_39),.co(co9_39),.a(pp10_30),.b(sum8_40),.ci(co8_39));
  fa u_csa9_40 (.s(sum9_40),.co(co9_40),.a(pp10_31),.b(sum8_41),.ci(co8_40));
  fa u_csa9_41 (.s(sum9_41),.co(co9_41),.a(pp10_32),.b(sum8_42),.ci(co8_41));
  fa u_csa9_42 (.s(sum9_42),.co(co9_42),.a(pp10_33),.b(sum8_43),.ci(co8_42));
  fa u_csa9_43 (.s(sum9_43),.co(co9_43),.a(pp10_34),.b(sum8_44),.ci(co8_43));
  assign sum9_44=pp10_35;
  assign co9_44=sig0;
  assign sum9_45=pp10_36;
  //CSA Row 10 
  ha u_csa10_0 (.s(sum10_0),.co(co10_0),.a(sum9_1),.b(co9_0));
  ha u_csa10_1 (.s(sum10_1),.co(co10_1),.a(sum9_2),.b(co9_1));
  ha u_csa10_2 (.s(sum10_2),.co(co10_2),.a(sum9_3),.b(co9_2));
  ha u_csa10_3 (.s(sum10_3),.co(co10_3),.a(sum9_4),.b(co9_3));
  ha u_csa10_4 (.s(sum10_4),.co(co10_4),.a(sum9_5),.b(co9_4));
  ha u_csa10_5 (.s(sum10_5),.co(co10_5),.a(sum9_6),.b(co9_5));
  ha u_csa10_6 (.s(sum10_6),.co(co10_6),.a(sum9_7),.b(co9_6));
  ha u_csa10_7 (.s(sum10_7),.co(co10_7),.a(sum9_8),.b(co9_7));
  ha u_csa10_8 (.s(sum10_8),.co(co10_8),.a(sum9_9),.b(co9_8));
  ha u_csa10_9 (.s(sum10_9),.co(co10_9),.a(sum9_10),.b(co9_9));
  fa u_csa10_10 (.s(sum10_10),.co(co10_10),.a(pp11_0),.b(sum9_11),.ci(co9_10));
  fa u_csa10_11 (.s(sum10_11),.co(co10_11),.a(pp11_1),.b(sum9_12),.ci(co9_11));
  fa u_csa10_12 (.s(sum10_12),.co(co10_12),.a(pp11_2),.b(sum9_13),.ci(co9_12));
  fa u_csa10_13 (.s(sum10_13),.co(co10_13),.a(pp11_3),.b(sum9_14),.ci(co9_13));
  fa u_csa10_14 (.s(sum10_14),.co(co10_14),.a(pp11_4),.b(sum9_15),.ci(co9_14));
  fa u_csa10_15 (.s(sum10_15),.co(co10_15),.a(pp11_5),.b(sum9_16),.ci(co9_15));
  fa u_csa10_16 (.s(sum10_16),.co(co10_16),.a(pp11_6),.b(sum9_17),.ci(co9_16));
  fa u_csa10_17 (.s(sum10_17),.co(co10_17),.a(pp11_7),.b(sum9_18),.ci(co9_17));
  fa u_csa10_18 (.s(sum10_18),.co(co10_18),.a(pp11_8),.b(sum9_19),.ci(co9_18));
  fa u_csa10_19 (.s(sum10_19),.co(co10_19),.a(pp11_9),.b(sum9_20),.ci(co9_19));
  fa u_csa10_20 (.s(sum10_20),.co(co10_20),.a(pp11_10),.b(sum9_21),.ci(co9_20));
  fa u_csa10_21 (.s(sum10_21),.co(co10_21),.a(pp11_11),.b(sum9_22),.ci(co9_21));
  fa u_csa10_22 (.s(sum10_22),.co(co10_22),.a(pp11_12),.b(sum9_23),.ci(co9_22));
  fa u_csa10_23 (.s(sum10_23),.co(co10_23),.a(pp11_13),.b(sum9_24),.ci(co9_23));
  fa u_csa10_24 (.s(sum10_24),.co(co10_24),.a(pp11_14),.b(sum9_25),.ci(co9_24));
  fa u_csa10_25 (.s(sum10_25),.co(co10_25),.a(pp11_15),.b(sum9_26),.ci(co9_25));
  fa u_csa10_26 (.s(sum10_26),.co(co10_26),.a(pp11_16),.b(sum9_27),.ci(co9_26));
  fa u_csa10_27 (.s(sum10_27),.co(co10_27),.a(pp11_17),.b(sum9_28),.ci(co9_27));
  fa u_csa10_28 (.s(sum10_28),.co(co10_28),.a(pp11_18),.b(sum9_29),.ci(co9_28));
  fa u_csa10_29 (.s(sum10_29),.co(co10_29),.a(pp11_19),.b(sum9_30),.ci(co9_29));
  fa u_csa10_30 (.s(sum10_30),.co(co10_30),.a(pp11_20),.b(sum9_31),.ci(co9_30));
  fa u_csa10_31 (.s(sum10_31),.co(co10_31),.a(pp11_21),.b(sum9_32),.ci(co9_31));
  fa u_csa10_32 (.s(sum10_32),.co(co10_32),.a(pp11_22),.b(sum9_33),.ci(co9_32));
  fa u_csa10_33 (.s(sum10_33),.co(co10_33),.a(pp11_23),.b(sum9_34),.ci(co9_33));
  fa u_csa10_34 (.s(sum10_34),.co(co10_34),.a(pp11_24),.b(sum9_35),.ci(co9_34));
  fa u_csa10_35 (.s(sum10_35),.co(co10_35),.a(pp11_25),.b(sum9_36),.ci(co9_35));
  fa u_csa10_36 (.s(sum10_36),.co(co10_36),.a(pp11_26),.b(sum9_37),.ci(co9_36));
  fa u_csa10_37 (.s(sum10_37),.co(co10_37),.a(pp11_27),.b(sum9_38),.ci(co9_37));
  fa u_csa10_38 (.s(sum10_38),.co(co10_38),.a(pp11_28),.b(sum9_39),.ci(co9_38));
  fa u_csa10_39 (.s(sum10_39),.co(co10_39),.a(pp11_29),.b(sum9_40),.ci(co9_39));
  fa u_csa10_40 (.s(sum10_40),.co(co10_40),.a(pp11_30),.b(sum9_41),.ci(co9_40));
  fa u_csa10_41 (.s(sum10_41),.co(co10_41),.a(pp11_31),.b(sum9_42),.ci(co9_41));
  fa u_csa10_42 (.s(sum10_42),.co(co10_42),.a(pp11_32),.b(sum9_43),.ci(co9_42));
  fa u_csa10_43 (.s(sum10_43),.co(co10_43),.a(pp11_33),.b(sum9_44),.ci(co9_43));
  fa u_csa10_44 (.s(sum10_44),.co(co10_44),.a(pp11_34),.b(sum9_45),.ci(co9_44));
  assign sum10_45=pp11_35;
  assign co10_45=sig0;
  assign sum10_46=pp11_36;
  //CSA Row 11 
  ha u_csa11_0 (.s(sum11_0),.co(co11_0),.a(sum10_1),.b(co10_0));
  ha u_csa11_1 (.s(sum11_1),.co(co11_1),.a(sum10_2),.b(co10_1));
  ha u_csa11_2 (.s(sum11_2),.co(co11_2),.a(sum10_3),.b(co10_2));
  ha u_csa11_3 (.s(sum11_3),.co(co11_3),.a(sum10_4),.b(co10_3));
  ha u_csa11_4 (.s(sum11_4),.co(co11_4),.a(sum10_5),.b(co10_4));
  ha u_csa11_5 (.s(sum11_5),.co(co11_5),.a(sum10_6),.b(co10_5));
  ha u_csa11_6 (.s(sum11_6),.co(co11_6),.a(sum10_7),.b(co10_6));
  ha u_csa11_7 (.s(sum11_7),.co(co11_7),.a(sum10_8),.b(co10_7));
  ha u_csa11_8 (.s(sum11_8),.co(co11_8),.a(sum10_9),.b(co10_8));
  ha u_csa11_9 (.s(sum11_9),.co(co11_9),.a(sum10_10),.b(co10_9));
  ha u_csa11_10 (.s(sum11_10),.co(co11_10),.a(sum10_11),.b(co10_10));
  fa u_csa11_11 (.s(sum11_11),.co(co11_11),.a(pp12_0),.b(sum10_12),.ci(co10_11));
  fa u_csa11_12 (.s(sum11_12),.co(co11_12),.a(pp12_1),.b(sum10_13),.ci(co10_12));
  fa u_csa11_13 (.s(sum11_13),.co(co11_13),.a(pp12_2),.b(sum10_14),.ci(co10_13));
  fa u_csa11_14 (.s(sum11_14),.co(co11_14),.a(pp12_3),.b(sum10_15),.ci(co10_14));
  fa u_csa11_15 (.s(sum11_15),.co(co11_15),.a(pp12_4),.b(sum10_16),.ci(co10_15));
  fa u_csa11_16 (.s(sum11_16),.co(co11_16),.a(pp12_5),.b(sum10_17),.ci(co10_16));
  fa u_csa11_17 (.s(sum11_17),.co(co11_17),.a(pp12_6),.b(sum10_18),.ci(co10_17));
  fa u_csa11_18 (.s(sum11_18),.co(co11_18),.a(pp12_7),.b(sum10_19),.ci(co10_18));
  fa u_csa11_19 (.s(sum11_19),.co(co11_19),.a(pp12_8),.b(sum10_20),.ci(co10_19));
  fa u_csa11_20 (.s(sum11_20),.co(co11_20),.a(pp12_9),.b(sum10_21),.ci(co10_20));
  fa u_csa11_21 (.s(sum11_21),.co(co11_21),.a(pp12_10),.b(sum10_22),.ci(co10_21));
  fa u_csa11_22 (.s(sum11_22),.co(co11_22),.a(pp12_11),.b(sum10_23),.ci(co10_22));
  fa u_csa11_23 (.s(sum11_23),.co(co11_23),.a(pp12_12),.b(sum10_24),.ci(co10_23));
  fa u_csa11_24 (.s(sum11_24),.co(co11_24),.a(pp12_13),.b(sum10_25),.ci(co10_24));
  fa u_csa11_25 (.s(sum11_25),.co(co11_25),.a(pp12_14),.b(sum10_26),.ci(co10_25));
  fa u_csa11_26 (.s(sum11_26),.co(co11_26),.a(pp12_15),.b(sum10_27),.ci(co10_26));
  fa u_csa11_27 (.s(sum11_27),.co(co11_27),.a(pp12_16),.b(sum10_28),.ci(co10_27));
  fa u_csa11_28 (.s(sum11_28),.co(co11_28),.a(pp12_17),.b(sum10_29),.ci(co10_28));
  fa u_csa11_29 (.s(sum11_29),.co(co11_29),.a(pp12_18),.b(sum10_30),.ci(co10_29));
  fa u_csa11_30 (.s(sum11_30),.co(co11_30),.a(pp12_19),.b(sum10_31),.ci(co10_30));
  fa u_csa11_31 (.s(sum11_31),.co(co11_31),.a(pp12_20),.b(sum10_32),.ci(co10_31));
  fa u_csa11_32 (.s(sum11_32),.co(co11_32),.a(pp12_21),.b(sum10_33),.ci(co10_32));
  fa u_csa11_33 (.s(sum11_33),.co(co11_33),.a(pp12_22),.b(sum10_34),.ci(co10_33));
  fa u_csa11_34 (.s(sum11_34),.co(co11_34),.a(pp12_23),.b(sum10_35),.ci(co10_34));
  fa u_csa11_35 (.s(sum11_35),.co(co11_35),.a(pp12_24),.b(sum10_36),.ci(co10_35));
  fa u_csa11_36 (.s(sum11_36),.co(co11_36),.a(pp12_25),.b(sum10_37),.ci(co10_36));
  fa u_csa11_37 (.s(sum11_37),.co(co11_37),.a(pp12_26),.b(sum10_38),.ci(co10_37));
  fa u_csa11_38 (.s(sum11_38),.co(co11_38),.a(pp12_27),.b(sum10_39),.ci(co10_38));
  fa u_csa11_39 (.s(sum11_39),.co(co11_39),.a(pp12_28),.b(sum10_40),.ci(co10_39));
  fa u_csa11_40 (.s(sum11_40),.co(co11_40),.a(pp12_29),.b(sum10_41),.ci(co10_40));
  fa u_csa11_41 (.s(sum11_41),.co(co11_41),.a(pp12_30),.b(sum10_42),.ci(co10_41));
  fa u_csa11_42 (.s(sum11_42),.co(co11_42),.a(pp12_31),.b(sum10_43),.ci(co10_42));
  fa u_csa11_43 (.s(sum11_43),.co(co11_43),.a(pp12_32),.b(sum10_44),.ci(co10_43));
  fa u_csa11_44 (.s(sum11_44),.co(co11_44),.a(pp12_33),.b(sum10_45),.ci(co10_44));
  fa u_csa11_45 (.s(sum11_45),.co(co11_45),.a(pp12_34),.b(sum10_46),.ci(co10_45));
  assign sum11_46=pp12_35;
  assign co11_46=sig0;
  assign sum11_47=pp12_36;
  //CSA Row 12 
  ha u_csa12_0 (.s(sum12_0),.co(co12_0),.a(sum11_1),.b(co11_0));
  ha u_csa12_1 (.s(sum12_1),.co(co12_1),.a(sum11_2),.b(co11_1));
  ha u_csa12_2 (.s(sum12_2),.co(co12_2),.a(sum11_3),.b(co11_2));
  ha u_csa12_3 (.s(sum12_3),.co(co12_3),.a(sum11_4),.b(co11_3));
  ha u_csa12_4 (.s(sum12_4),.co(co12_4),.a(sum11_5),.b(co11_4));
  ha u_csa12_5 (.s(sum12_5),.co(co12_5),.a(sum11_6),.b(co11_5));
  ha u_csa12_6 (.s(sum12_6),.co(co12_6),.a(sum11_7),.b(co11_6));
  ha u_csa12_7 (.s(sum12_7),.co(co12_7),.a(sum11_8),.b(co11_7));
  ha u_csa12_8 (.s(sum12_8),.co(co12_8),.a(sum11_9),.b(co11_8));
  ha u_csa12_9 (.s(sum12_9),.co(co12_9),.a(sum11_10),.b(co11_9));
  ha u_csa12_10 (.s(sum12_10),.co(co12_10),.a(sum11_11),.b(co11_10));
  ha u_csa12_11 (.s(sum12_11),.co(co12_11),.a(sum11_12),.b(co11_11));
  fa u_csa12_12 (.s(sum12_12),.co(co12_12),.a(pp13_0),.b(sum11_13),.ci(co11_12));
  fa u_csa12_13 (.s(sum12_13),.co(co12_13),.a(pp13_1),.b(sum11_14),.ci(co11_13));
  fa u_csa12_14 (.s(sum12_14),.co(co12_14),.a(pp13_2),.b(sum11_15),.ci(co11_14));
  fa u_csa12_15 (.s(sum12_15),.co(co12_15),.a(pp13_3),.b(sum11_16),.ci(co11_15));
  fa u_csa12_16 (.s(sum12_16),.co(co12_16),.a(pp13_4),.b(sum11_17),.ci(co11_16));
  fa u_csa12_17 (.s(sum12_17),.co(co12_17),.a(pp13_5),.b(sum11_18),.ci(co11_17));
  fa u_csa12_18 (.s(sum12_18),.co(co12_18),.a(pp13_6),.b(sum11_19),.ci(co11_18));
  fa u_csa12_19 (.s(sum12_19),.co(co12_19),.a(pp13_7),.b(sum11_20),.ci(co11_19));
  fa u_csa12_20 (.s(sum12_20),.co(co12_20),.a(pp13_8),.b(sum11_21),.ci(co11_20));
  fa u_csa12_21 (.s(sum12_21),.co(co12_21),.a(pp13_9),.b(sum11_22),.ci(co11_21));
  fa u_csa12_22 (.s(sum12_22),.co(co12_22),.a(pp13_10),.b(sum11_23),.ci(co11_22));
  fa u_csa12_23 (.s(sum12_23),.co(co12_23),.a(pp13_11),.b(sum11_24),.ci(co11_23));
  fa u_csa12_24 (.s(sum12_24),.co(co12_24),.a(pp13_12),.b(sum11_25),.ci(co11_24));
  fa u_csa12_25 (.s(sum12_25),.co(co12_25),.a(pp13_13),.b(sum11_26),.ci(co11_25));
  fa u_csa12_26 (.s(sum12_26),.co(co12_26),.a(pp13_14),.b(sum11_27),.ci(co11_26));
  fa u_csa12_27 (.s(sum12_27),.co(co12_27),.a(pp13_15),.b(sum11_28),.ci(co11_27));
  fa u_csa12_28 (.s(sum12_28),.co(co12_28),.a(pp13_16),.b(sum11_29),.ci(co11_28));
  fa u_csa12_29 (.s(sum12_29),.co(co12_29),.a(pp13_17),.b(sum11_30),.ci(co11_29));
  fa u_csa12_30 (.s(sum12_30),.co(co12_30),.a(pp13_18),.b(sum11_31),.ci(co11_30));
  fa u_csa12_31 (.s(sum12_31),.co(co12_31),.a(pp13_19),.b(sum11_32),.ci(co11_31));
  fa u_csa12_32 (.s(sum12_32),.co(co12_32),.a(pp13_20),.b(sum11_33),.ci(co11_32));
  fa u_csa12_33 (.s(sum12_33),.co(co12_33),.a(pp13_21),.b(sum11_34),.ci(co11_33));
  fa u_csa12_34 (.s(sum12_34),.co(co12_34),.a(pp13_22),.b(sum11_35),.ci(co11_34));
  fa u_csa12_35 (.s(sum12_35),.co(co12_35),.a(pp13_23),.b(sum11_36),.ci(co11_35));
  fa u_csa12_36 (.s(sum12_36),.co(co12_36),.a(pp13_24),.b(sum11_37),.ci(co11_36));
  fa u_csa12_37 (.s(sum12_37),.co(co12_37),.a(pp13_25),.b(sum11_38),.ci(co11_37));
  fa u_csa12_38 (.s(sum12_38),.co(co12_38),.a(pp13_26),.b(sum11_39),.ci(co11_38));
  fa u_csa12_39 (.s(sum12_39),.co(co12_39),.a(pp13_27),.b(sum11_40),.ci(co11_39));
  fa u_csa12_40 (.s(sum12_40),.co(co12_40),.a(pp13_28),.b(sum11_41),.ci(co11_40));
  fa u_csa12_41 (.s(sum12_41),.co(co12_41),.a(pp13_29),.b(sum11_42),.ci(co11_41));
  fa u_csa12_42 (.s(sum12_42),.co(co12_42),.a(pp13_30),.b(sum11_43),.ci(co11_42));
  fa u_csa12_43 (.s(sum12_43),.co(co12_43),.a(pp13_31),.b(sum11_44),.ci(co11_43));
  fa u_csa12_44 (.s(sum12_44),.co(co12_44),.a(pp13_32),.b(sum11_45),.ci(co11_44));
  fa u_csa12_45 (.s(sum12_45),.co(co12_45),.a(pp13_33),.b(sum11_46),.ci(co11_45));
  fa u_csa12_46 (.s(sum12_46),.co(co12_46),.a(pp13_34),.b(sum11_47),.ci(co11_46));
  assign sum12_47=pp13_35;
  assign co12_47=sig0;
  assign sum12_48=pp13_36;
  //CSA Row 13 
  ha u_csa13_0 (.s(sum13_0),.co(co13_0),.a(sum12_1),.b(co12_0));
  ha u_csa13_1 (.s(sum13_1),.co(co13_1),.a(sum12_2),.b(co12_1));
  ha u_csa13_2 (.s(sum13_2),.co(co13_2),.a(sum12_3),.b(co12_2));
  ha u_csa13_3 (.s(sum13_3),.co(co13_3),.a(sum12_4),.b(co12_3));
  ha u_csa13_4 (.s(sum13_4),.co(co13_4),.a(sum12_5),.b(co12_4));
  ha u_csa13_5 (.s(sum13_5),.co(co13_5),.a(sum12_6),.b(co12_5));
  ha u_csa13_6 (.s(sum13_6),.co(co13_6),.a(sum12_7),.b(co12_6));
  ha u_csa13_7 (.s(sum13_7),.co(co13_7),.a(sum12_8),.b(co12_7));
  ha u_csa13_8 (.s(sum13_8),.co(co13_8),.a(sum12_9),.b(co12_8));
  ha u_csa13_9 (.s(sum13_9),.co(co13_9),.a(sum12_10),.b(co12_9));
  ha u_csa13_10 (.s(sum13_10),.co(co13_10),.a(sum12_11),.b(co12_10));
  ha u_csa13_11 (.s(sum13_11),.co(co13_11),.a(sum12_12),.b(co12_11));
  ha u_csa13_12 (.s(sum13_12),.co(co13_12),.a(sum12_13),.b(co12_12));
  fa u_csa13_13 (.s(sum13_13),.co(co13_13),.a(pp14_0),.b(sum12_14),.ci(co12_13));
  fa u_csa13_14 (.s(sum13_14),.co(co13_14),.a(pp14_1),.b(sum12_15),.ci(co12_14));
  fa u_csa13_15 (.s(sum13_15),.co(co13_15),.a(pp14_2),.b(sum12_16),.ci(co12_15));
  fa u_csa13_16 (.s(sum13_16),.co(co13_16),.a(pp14_3),.b(sum12_17),.ci(co12_16));
  fa u_csa13_17 (.s(sum13_17),.co(co13_17),.a(pp14_4),.b(sum12_18),.ci(co12_17));
  fa u_csa13_18 (.s(sum13_18),.co(co13_18),.a(pp14_5),.b(sum12_19),.ci(co12_18));
  fa u_csa13_19 (.s(sum13_19),.co(co13_19),.a(pp14_6),.b(sum12_20),.ci(co12_19));
  fa u_csa13_20 (.s(sum13_20),.co(co13_20),.a(pp14_7),.b(sum12_21),.ci(co12_20));
  fa u_csa13_21 (.s(sum13_21),.co(co13_21),.a(pp14_8),.b(sum12_22),.ci(co12_21));
  fa u_csa13_22 (.s(sum13_22),.co(co13_22),.a(pp14_9),.b(sum12_23),.ci(co12_22));
  fa u_csa13_23 (.s(sum13_23),.co(co13_23),.a(pp14_10),.b(sum12_24),.ci(co12_23));
  fa u_csa13_24 (.s(sum13_24),.co(co13_24),.a(pp14_11),.b(sum12_25),.ci(co12_24));
  fa u_csa13_25 (.s(sum13_25),.co(co13_25),.a(pp14_12),.b(sum12_26),.ci(co12_25));
  fa u_csa13_26 (.s(sum13_26),.co(co13_26),.a(pp14_13),.b(sum12_27),.ci(co12_26));
  fa u_csa13_27 (.s(sum13_27),.co(co13_27),.a(pp14_14),.b(sum12_28),.ci(co12_27));
  fa u_csa13_28 (.s(sum13_28),.co(co13_28),.a(pp14_15),.b(sum12_29),.ci(co12_28));
  fa u_csa13_29 (.s(sum13_29),.co(co13_29),.a(pp14_16),.b(sum12_30),.ci(co12_29));
  fa u_csa13_30 (.s(sum13_30),.co(co13_30),.a(pp14_17),.b(sum12_31),.ci(co12_30));
  fa u_csa13_31 (.s(sum13_31),.co(co13_31),.a(pp14_18),.b(sum12_32),.ci(co12_31));
  fa u_csa13_32 (.s(sum13_32),.co(co13_32),.a(pp14_19),.b(sum12_33),.ci(co12_32));
  fa u_csa13_33 (.s(sum13_33),.co(co13_33),.a(pp14_20),.b(sum12_34),.ci(co12_33));
  fa u_csa13_34 (.s(sum13_34),.co(co13_34),.a(pp14_21),.b(sum12_35),.ci(co12_34));
  fa u_csa13_35 (.s(sum13_35),.co(co13_35),.a(pp14_22),.b(sum12_36),.ci(co12_35));
  fa u_csa13_36 (.s(sum13_36),.co(co13_36),.a(pp14_23),.b(sum12_37),.ci(co12_36));
  fa u_csa13_37 (.s(sum13_37),.co(co13_37),.a(pp14_24),.b(sum12_38),.ci(co12_37));
  fa u_csa13_38 (.s(sum13_38),.co(co13_38),.a(pp14_25),.b(sum12_39),.ci(co12_38));
  fa u_csa13_39 (.s(sum13_39),.co(co13_39),.a(pp14_26),.b(sum12_40),.ci(co12_39));
  fa u_csa13_40 (.s(sum13_40),.co(co13_40),.a(pp14_27),.b(sum12_41),.ci(co12_40));
  fa u_csa13_41 (.s(sum13_41),.co(co13_41),.a(pp14_28),.b(sum12_42),.ci(co12_41));
  fa u_csa13_42 (.s(sum13_42),.co(co13_42),.a(pp14_29),.b(sum12_43),.ci(co12_42));
  fa u_csa13_43 (.s(sum13_43),.co(co13_43),.a(pp14_30),.b(sum12_44),.ci(co12_43));
  fa u_csa13_44 (.s(sum13_44),.co(co13_44),.a(pp14_31),.b(sum12_45),.ci(co12_44));
  fa u_csa13_45 (.s(sum13_45),.co(co13_45),.a(pp14_32),.b(sum12_46),.ci(co12_45));
  fa u_csa13_46 (.s(sum13_46),.co(co13_46),.a(pp14_33),.b(sum12_47),.ci(co12_46));
  fa u_csa13_47 (.s(sum13_47),.co(co13_47),.a(pp14_34),.b(sum12_48),.ci(co12_47));
  assign sum13_48=pp14_35;
  assign co13_48=sig0;
  assign sum13_49=pp14_36;
  //CSA Row 14 
  ha u_csa14_0 (.s(sum14_0),.co(co14_0),.a(sum13_1),.b(co13_0));
  ha u_csa14_1 (.s(sum14_1),.co(co14_1),.a(sum13_2),.b(co13_1));
  ha u_csa14_2 (.s(sum14_2),.co(co14_2),.a(sum13_3),.b(co13_2));
  ha u_csa14_3 (.s(sum14_3),.co(co14_3),.a(sum13_4),.b(co13_3));
  ha u_csa14_4 (.s(sum14_4),.co(co14_4),.a(sum13_5),.b(co13_4));
  ha u_csa14_5 (.s(sum14_5),.co(co14_5),.a(sum13_6),.b(co13_5));
  ha u_csa14_6 (.s(sum14_6),.co(co14_6),.a(sum13_7),.b(co13_6));
  ha u_csa14_7 (.s(sum14_7),.co(co14_7),.a(sum13_8),.b(co13_7));
  ha u_csa14_8 (.s(sum14_8),.co(co14_8),.a(sum13_9),.b(co13_8));
  ha u_csa14_9 (.s(sum14_9),.co(co14_9),.a(sum13_10),.b(co13_9));
  ha u_csa14_10 (.s(sum14_10),.co(co14_10),.a(sum13_11),.b(co13_10));
  ha u_csa14_11 (.s(sum14_11),.co(co14_11),.a(sum13_12),.b(co13_11));
  ha u_csa14_12 (.s(sum14_12),.co(co14_12),.a(sum13_13),.b(co13_12));
  ha u_csa14_13 (.s(sum14_13),.co(co14_13),.a(sum13_14),.b(co13_13));
  fa u_csa14_14 (.s(sum14_14),.co(co14_14),.a(pp15_0),.b(sum13_15),.ci(co13_14));
  fa u_csa14_15 (.s(sum14_15),.co(co14_15),.a(pp15_1),.b(sum13_16),.ci(co13_15));
  fa u_csa14_16 (.s(sum14_16),.co(co14_16),.a(pp15_2),.b(sum13_17),.ci(co13_16));
  fa u_csa14_17 (.s(sum14_17),.co(co14_17),.a(pp15_3),.b(sum13_18),.ci(co13_17));
  fa u_csa14_18 (.s(sum14_18),.co(co14_18),.a(pp15_4),.b(sum13_19),.ci(co13_18));
  fa u_csa14_19 (.s(sum14_19),.co(co14_19),.a(pp15_5),.b(sum13_20),.ci(co13_19));
  fa u_csa14_20 (.s(sum14_20),.co(co14_20),.a(pp15_6),.b(sum13_21),.ci(co13_20));
  fa u_csa14_21 (.s(sum14_21),.co(co14_21),.a(pp15_7),.b(sum13_22),.ci(co13_21));
  fa u_csa14_22 (.s(sum14_22),.co(co14_22),.a(pp15_8),.b(sum13_23),.ci(co13_22));
  fa u_csa14_23 (.s(sum14_23),.co(co14_23),.a(pp15_9),.b(sum13_24),.ci(co13_23));
  fa u_csa14_24 (.s(sum14_24),.co(co14_24),.a(pp15_10),.b(sum13_25),.ci(co13_24));
  fa u_csa14_25 (.s(sum14_25),.co(co14_25),.a(pp15_11),.b(sum13_26),.ci(co13_25));
  fa u_csa14_26 (.s(sum14_26),.co(co14_26),.a(pp15_12),.b(sum13_27),.ci(co13_26));
  fa u_csa14_27 (.s(sum14_27),.co(co14_27),.a(pp15_13),.b(sum13_28),.ci(co13_27));
  fa u_csa14_28 (.s(sum14_28),.co(co14_28),.a(pp15_14),.b(sum13_29),.ci(co13_28));
  fa u_csa14_29 (.s(sum14_29),.co(co14_29),.a(pp15_15),.b(sum13_30),.ci(co13_29));
  fa u_csa14_30 (.s(sum14_30),.co(co14_30),.a(pp15_16),.b(sum13_31),.ci(co13_30));
  fa u_csa14_31 (.s(sum14_31),.co(co14_31),.a(pp15_17),.b(sum13_32),.ci(co13_31));
  fa u_csa14_32 (.s(sum14_32),.co(co14_32),.a(pp15_18),.b(sum13_33),.ci(co13_32));
  fa u_csa14_33 (.s(sum14_33),.co(co14_33),.a(pp15_19),.b(sum13_34),.ci(co13_33));
  fa u_csa14_34 (.s(sum14_34),.co(co14_34),.a(pp15_20),.b(sum13_35),.ci(co13_34));
  fa u_csa14_35 (.s(sum14_35),.co(co14_35),.a(pp15_21),.b(sum13_36),.ci(co13_35));
  fa u_csa14_36 (.s(sum14_36),.co(co14_36),.a(pp15_22),.b(sum13_37),.ci(co13_36));
  fa u_csa14_37 (.s(sum14_37),.co(co14_37),.a(pp15_23),.b(sum13_38),.ci(co13_37));
  fa u_csa14_38 (.s(sum14_38),.co(co14_38),.a(pp15_24),.b(sum13_39),.ci(co13_38));
  fa u_csa14_39 (.s(sum14_39),.co(co14_39),.a(pp15_25),.b(sum13_40),.ci(co13_39));
  fa u_csa14_40 (.s(sum14_40),.co(co14_40),.a(pp15_26),.b(sum13_41),.ci(co13_40));
  fa u_csa14_41 (.s(sum14_41),.co(co14_41),.a(pp15_27),.b(sum13_42),.ci(co13_41));
  fa u_csa14_42 (.s(sum14_42),.co(co14_42),.a(pp15_28),.b(sum13_43),.ci(co13_42));
  fa u_csa14_43 (.s(sum14_43),.co(co14_43),.a(pp15_29),.b(sum13_44),.ci(co13_43));
  fa u_csa14_44 (.s(sum14_44),.co(co14_44),.a(pp15_30),.b(sum13_45),.ci(co13_44));
  fa u_csa14_45 (.s(sum14_45),.co(co14_45),.a(pp15_31),.b(sum13_46),.ci(co13_45));
  fa u_csa14_46 (.s(sum14_46),.co(co14_46),.a(pp15_32),.b(sum13_47),.ci(co13_46));
  fa u_csa14_47 (.s(sum14_47),.co(co14_47),.a(pp15_33),.b(sum13_48),.ci(co13_47));
  fa u_csa14_48 (.s(sum14_48),.co(co14_48),.a(pp15_34),.b(sum13_49),.ci(co13_48));
  assign sum14_49=pp15_35;
  assign co14_49=sig0;
  //CSA Row 15 
  ha u_csa15_0 (.s(sum15_0),.co(co15_0),.a(sum14_1),.b(co14_0));
  ha u_csa15_1 (.s(sum15_1),.co(co15_1),.a(sum14_2),.b(co14_1));
  ha u_csa15_2 (.s(sum15_2),.co(co15_2),.a(sum14_3),.b(co14_2));
  ha u_csa15_3 (.s(sum15_3),.co(co15_3),.a(sum14_4),.b(co14_3));
  ha u_csa15_4 (.s(sum15_4),.co(co15_4),.a(sum14_5),.b(co14_4));
  ha u_csa15_5 (.s(sum15_5),.co(co15_5),.a(sum14_6),.b(co14_5));
  ha u_csa15_6 (.s(sum15_6),.co(co15_6),.a(sum14_7),.b(co14_6));
  ha u_csa15_7 (.s(sum15_7),.co(co15_7),.a(sum14_8),.b(co14_7));
  ha u_csa15_8 (.s(sum15_8),.co(co15_8),.a(sum14_9),.b(co14_8));
  ha u_csa15_9 (.s(sum15_9),.co(co15_9),.a(sum14_10),.b(co14_9));
  ha u_csa15_10 (.s(sum15_10),.co(co15_10),.a(sum14_11),.b(co14_10));
  ha u_csa15_11 (.s(sum15_11),.co(co15_11),.a(sum14_12),.b(co14_11));
  ha u_csa15_12 (.s(sum15_12),.co(co15_12),.a(sum14_13),.b(co14_12));
  ha u_csa15_13 (.s(sum15_13),.co(co15_13),.a(sum14_14),.b(co14_13));
  ha u_csa15_14 (.s(sum15_14),.co(co15_14),.a(sum14_15),.b(co14_14));
  fa u_csa15_15 (.s(sum15_15),.co(co15_15),.a(pp16_0),.b(sum14_16),.ci(co14_15));
  fa u_csa15_16 (.s(sum15_16),.co(co15_16),.a(pp16_1),.b(sum14_17),.ci(co14_16));
  fa u_csa15_17 (.s(sum15_17),.co(co15_17),.a(pp16_2),.b(sum14_18),.ci(co14_17));
  fa u_csa15_18 (.s(sum15_18),.co(co15_18),.a(pp16_3),.b(sum14_19),.ci(co14_18));
  fa u_csa15_19 (.s(sum15_19),.co(co15_19),.a(pp16_4),.b(sum14_20),.ci(co14_19));
  fa u_csa15_20 (.s(sum15_20),.co(co15_20),.a(pp16_5),.b(sum14_21),.ci(co14_20));
  fa u_csa15_21 (.s(sum15_21),.co(co15_21),.a(pp16_6),.b(sum14_22),.ci(co14_21));
  fa u_csa15_22 (.s(sum15_22),.co(co15_22),.a(pp16_7),.b(sum14_23),.ci(co14_22));
  fa u_csa15_23 (.s(sum15_23),.co(co15_23),.a(pp16_8),.b(sum14_24),.ci(co14_23));
  fa u_csa15_24 (.s(sum15_24),.co(co15_24),.a(pp16_9),.b(sum14_25),.ci(co14_24));
  fa u_csa15_25 (.s(sum15_25),.co(co15_25),.a(pp16_10),.b(sum14_26),.ci(co14_25));
  fa u_csa15_26 (.s(sum15_26),.co(co15_26),.a(pp16_11),.b(sum14_27),.ci(co14_26));
  fa u_csa15_27 (.s(sum15_27),.co(co15_27),.a(pp16_12),.b(sum14_28),.ci(co14_27));
  fa u_csa15_28 (.s(sum15_28),.co(co15_28),.a(pp16_13),.b(sum14_29),.ci(co14_28));
  fa u_csa15_29 (.s(sum15_29),.co(co15_29),.a(pp16_14),.b(sum14_30),.ci(co14_29));
  fa u_csa15_30 (.s(sum15_30),.co(co15_30),.a(pp16_15),.b(sum14_31),.ci(co14_30));
  fa u_csa15_31 (.s(sum15_31),.co(co15_31),.a(pp16_16),.b(sum14_32),.ci(co14_31));
  fa u_csa15_32 (.s(sum15_32),.co(co15_32),.a(pp16_17),.b(sum14_33),.ci(co14_32));
  fa u_csa15_33 (.s(sum15_33),.co(co15_33),.a(pp16_18),.b(sum14_34),.ci(co14_33));
  fa u_csa15_34 (.s(sum15_34),.co(co15_34),.a(pp16_19),.b(sum14_35),.ci(co14_34));
  fa u_csa15_35 (.s(sum15_35),.co(co15_35),.a(pp16_20),.b(sum14_36),.ci(co14_35));
  fa u_csa15_36 (.s(sum15_36),.co(co15_36),.a(pp16_21),.b(sum14_37),.ci(co14_36));
  fa u_csa15_37 (.s(sum15_37),.co(co15_37),.a(pp16_22),.b(sum14_38),.ci(co14_37));
  fa u_csa15_38 (.s(sum15_38),.co(co15_38),.a(pp16_23),.b(sum14_39),.ci(co14_38));
  fa u_csa15_39 (.s(sum15_39),.co(co15_39),.a(pp16_24),.b(sum14_40),.ci(co14_39));
  fa u_csa15_40 (.s(sum15_40),.co(co15_40),.a(pp16_25),.b(sum14_41),.ci(co14_40));
  fa u_csa15_41 (.s(sum15_41),.co(co15_41),.a(pp16_26),.b(sum14_42),.ci(co14_41));
  fa u_csa15_42 (.s(sum15_42),.co(co15_42),.a(pp16_27),.b(sum14_43),.ci(co14_42));
  fa u_csa15_43 (.s(sum15_43),.co(co15_43),.a(pp16_28),.b(sum14_44),.ci(co14_43));
  fa u_csa15_44 (.s(sum15_44),.co(co15_44),.a(pp16_29),.b(sum14_45),.ci(co14_44));
  fa u_csa15_45 (.s(sum15_45),.co(co15_45),.a(pp16_30),.b(sum14_46),.ci(co14_45));
  fa u_csa15_46 (.s(sum15_46),.co(co15_46),.a(pp16_31),.b(sum14_47),.ci(co14_46));
  fa u_csa15_47 (.s(sum15_47),.co(co15_47),.a(pp16_32),.b(sum14_48),.ci(co14_47));
  fa u_csa15_48 (.s(sum15_48),.co(co15_48),.a(pp16_33),.b(sum14_49),.ci(co14_48));
  assign p[0]=sum0_0;
  assign p[1]=sum1_0;
  assign p[2]=sum2_0;
  assign p[3]=sum3_0;
  assign p[4]=sum4_0;
  assign p[5]=sum5_0;
  assign p[6]=sum6_0;
  assign p[7]=sum7_0;
  assign p[8]=sum8_0;
  assign p[9]=sum9_0;
  assign p[10]=sum10_0;
  assign p[11]=sum11_0;
  assign p[12]=sum12_0;
  assign p[13]=sum13_0;
  assign p[14]=sum14_0;
  assign p[15]=sum15_0;
  assign s_vec[0]=sum15_1;
  assign s_vec[1]=sum15_2;
  assign s_vec[2]=sum15_3;
  assign s_vec[3]=sum15_4;
  assign s_vec[4]=sum15_5;
  assign s_vec[5]=sum15_6;
  assign s_vec[6]=sum15_7;
  assign s_vec[7]=sum15_8;
  assign s_vec[8]=sum15_9;
  assign s_vec[9]=sum15_10;
  assign s_vec[10]=sum15_11;
  assign s_vec[11]=sum15_12;
  assign s_vec[12]=sum15_13;
  assign s_vec[13]=sum15_14;
  assign s_vec[14]=sum15_15;
  assign s_vec[15]=sum15_16;
  assign s_vec[16]=sum15_17;
  assign s_vec[17]=sum15_18;
  assign s_vec[18]=sum15_19;
  assign s_vec[19]=sum15_20;
  assign s_vec[20]=sum15_21;
  assign s_vec[21]=sum15_22;
  assign s_vec[22]=sum15_23;
  assign s_vec[23]=sum15_24;
  assign s_vec[24]=sum15_25;
  assign s_vec[25]=sum15_26;
  assign s_vec[26]=sum15_27;
  assign s_vec[27]=sum15_28;
  assign s_vec[28]=sum15_29;
  assign s_vec[29]=sum15_30;
  assign s_vec[30]=sum15_31;
  assign s_vec[31]=sum15_32;
  assign s_vec[32]=sum15_33;
  assign s_vec[33]=sum15_34;
  assign s_vec[34]=sum15_35;
  assign s_vec[35]=sum15_36;
  assign s_vec[36]=sum15_37;
  assign s_vec[37]=sum15_38;
  assign s_vec[38]=sum15_39;
  assign s_vec[39]=sum15_40;
  assign s_vec[40]=sum15_41;
  assign s_vec[41]=sum15_42;
  assign s_vec[42]=sum15_43;
  assign s_vec[43]=sum15_44;
  assign s_vec[44]=sum15_45;
  assign s_vec[45]=sum15_46;
  assign s_vec[46]=sum15_47;
  assign s_vec[47]=sum15_48;
  assign c_vec[0]=co15_0;
  assign c_vec[1]=co15_1;
  assign c_vec[2]=co15_2;
  assign c_vec[3]=co15_3;
  assign c_vec[4]=co15_4;
  assign c_vec[5]=co15_5;
  assign c_vec[6]=co15_6;
  assign c_vec[7]=co15_7;
  assign c_vec[8]=co15_8;
  assign c_vec[9]=co15_9;
  assign c_vec[10]=co15_10;
  assign c_vec[11]=co15_11;
  assign c_vec[12]=co15_12;
  assign c_vec[13]=co15_13;
  assign c_vec[14]=co15_14;
  assign c_vec[15]=co15_15;
  assign c_vec[16]=co15_16;
  assign c_vec[17]=co15_17;
  assign c_vec[18]=co15_18;
  assign c_vec[19]=co15_19;
  assign c_vec[20]=co15_20;
  assign c_vec[21]=co15_21;
  assign c_vec[22]=co15_22;
  assign c_vec[23]=co15_23;
  assign c_vec[24]=co15_24;
  assign c_vec[25]=co15_25;
  assign c_vec[26]=co15_26;
  assign c_vec[27]=co15_27;
  assign c_vec[28]=co15_28;
  assign c_vec[29]=co15_29;
  assign c_vec[30]=co15_30;
  assign c_vec[31]=co15_31;
  assign c_vec[32]=co15_32;
  assign c_vec[33]=co15_33;
  assign c_vec[34]=co15_34;
  assign c_vec[35]=co15_35;
  assign c_vec[36]=co15_36;
  assign c_vec[37]=co15_37;
  assign c_vec[38]=co15_38;
  assign c_vec[39]=co15_39;
  assign c_vec[40]=co15_40;
  assign c_vec[41]=co15_41;
  assign c_vec[42]=co15_42;
  assign c_vec[43]=co15_43;
  assign c_vec[44]=co15_44;
  assign c_vec[45]=co15_45;
  assign c_vec[46]=co15_46;
  assign c_vec[47]=co15_47;
  addripple_n #(.WIDTH(48))  u_add48 (.co(add_co),.s(p[63:16]),.a(s_vec),.b(c_vec));
 endmodule
